// Verilog simulation library for c35_IOLIB_ANA_3B_4M
// Owner: austriamicrosystems AG  HIT-Kit: Digital
module APRIO1K5P_3B (PAD,Z);
  inout PAD ;
  inout Z ;
endmodule
module APRIO200P_3B (PAD,Z);
  inout PAD ;
  inout Z ;
endmodule
module APRIO50P_3B (PAD,Z);
  inout PAD ;
  inout Z ;
endmodule
module APRIO500P_3B (PAD,Z);
  inout PAD ;
  inout Z ;
endmodule
module AVSUBP_3B (A);
  input A ;
endmodule
module APRIOWP_3B (PAD,Z);
  inout PAD ;
  inout Z ;
endmodule
module AGND3ALLP_3B (A);
  input A ;
endmodule
module AGND5ALLP_3B (A);
  input A ;
endmodule
module AVDD3ALLP_3B (A);
  input A ;
endmodule
module AVDD5ALLP_3B (A);
  input A ;
endmodule
module APRIOP_3B (PAD,Z);
  inout PAD ;
  inout Z ;
endmodule
module ARAILPROT3P_3B;
endmodule
module ARAILPRO5P_3B;
endmodule
