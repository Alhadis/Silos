// Verilog simulation library for c35_IOLIBC_ANA_3B_4M
// Owner: austriamicrosystems AG  HIT-Kit: Digital
module APRIO1K5C_3B (PAD,Z);
  inout PAD ;
  inout Z ;
endmodule
module APRIO200C_3B (PAD,Z);
  inout PAD ;
  inout Z ;
endmodule
module APRIO50C_3B (PAD,Z);
  inout PAD ;
  inout Z ;
endmodule
module APRIO500C_3B (PAD,Z);
  inout PAD ;
  inout Z ;
endmodule
module AVSUBC_3B (A);
  input A ;
endmodule
module APRIOWC1_3B (PAD,Z);
  inout PAD ;
  inout Z ;
endmodule
module AGND3ALLC_3B (A);
  input A ;
endmodule
module AGND5ALLC_3B (A);
  input A ;
endmodule
module AVDD3ALLC_3B (A);
  input A ;
endmodule
module AVDD5ALLC_3B (A);
  input A ;
endmodule
module APRIOC_3B (PAD,Z);
  inout PAD ;
  inout Z ;
endmodule
module ARAILPROT3C_3B;
endmodule
module ARAILPROT5C_3B;
endmodule
