
module system (
	clk_clk,
	reset_reset_n,
	rtc_module_0_conduit_end_export,
	rtc_module_0_conduit_end_1_export,
	rtc_module_0_conduit_end_2_export,
	rtc_module_0_conduit_end_3_export,
	rtc_module_0_conduit_end_4_export,
	rtc_module_0_conduit_end_5_export);	

	input		clk_clk;
	input		reset_reset_n;
	output	[3:0]	rtc_module_0_conduit_end_export;
	output		rtc_module_0_conduit_end_1_export;
	output	[7:0]	rtc_module_0_conduit_end_2_export;
	input	[7:0]	rtc_module_0_conduit_end_3_export;
	input	[3:0]	rtc_module_0_conduit_end_4_export;
	output	[5:0]	rtc_module_0_conduit_end_5_export;
endmodule
