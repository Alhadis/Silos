`timescale 1ns/100ps

module alu_shift_tb;

reg clock = 0;
integer dut_error = 0;

reg   [1:0] sfn;
reg  [31:0] a;
reg   [4:0] b;
wire [31:0] y;

// -------------------------------------------------------
// CLOCK GENERATION
// -------------------------------------------------------

always begin
	clock=0; #4;  // 125 MHz
	clock=1; #4;
end

// -------------------------------------------------------
// INITIALIZATION
// -------------------------------------------------------

initial begin
	if ($test$plusargs("vcd")) begin
		$dumpfile ("alu_shift_tb.vcd");
		$dumpvars (5, alu_shift_tb, dut);
	end
end

// -------------------------------------------------------
// TEST CASES
// -------------------------------------------------------

task test_case;
    input [38:0] inputs;
    input [31:0] expected_output;
	input integer line;
    begin
        {sfn, a, b} <= inputs;
        @(posedge clock)
        if (y == expected_output) begin
            $display("pass:  sfn=%01x, a=%08x, b=%02x => y=%08x",
                     inputs[38:37], inputs[36:5], inputs[4:0],
                     y);
        end else begin
            $display("FAIL:  sfn=%01x, a=%08x, b=%02x => y=%08x (expected %08x)",
                     inputs[38:37], inputs[36:5], inputs[4:0],
                     y,
                     expected_output);
			$error("");
			$display("       test_case at line %d", line);
			dut_error = dut_error + 1;
        end
    end
endtask

initial begin
    @(posedge clock);
    $display("");
	test_case({2'b00, 32'b00000000000000000000000000000000, 5'b00000}, 32'b00000000000000000000000000000000, `__LINE__); //   1: fn=SHL, a=0X00000000, b= 0, y=0X00000000
	test_case({2'b01, 32'b00000000000000000000000000000000, 5'b00000}, 32'b00000000000000000000000000000000, `__LINE__); //   2: fn=SHR, a=0X00000000, b= 0, y=0X00000000
	test_case({2'b11, 32'b00000000000000000000000000000000, 5'b00000}, 32'b00000000000000000000000000000000, `__LINE__); //   3: fn=SRA, a=0X00000000, b= 0, y=0X00000000
	test_case({2'b00, 32'b00000000000000000000000000000000, 5'b00001}, 32'b00000000000000000000000000000000, `__LINE__); //   4: fn=SHL, a=0X00000000, b= 1, y=0X00000000
	test_case({2'b01, 32'b00000000000000000000000000000000, 5'b00001}, 32'b00000000000000000000000000000000, `__LINE__); //   5: fn=SHR, a=0X00000000, b= 1, y=0X00000000
	test_case({2'b11, 32'b00000000000000000000000000000000, 5'b00001}, 32'b00000000000000000000000000000000, `__LINE__); //   6: fn=SRA, a=0X00000000, b= 1, y=0X00000000
	test_case({2'b00, 32'b00000000000000000000000000000000, 5'b00010}, 32'b00000000000000000000000000000000, `__LINE__); //   7: fn=SHL, a=0X00000000, b= 2, y=0X00000000
	test_case({2'b01, 32'b00000000000000000000000000000000, 5'b00010}, 32'b00000000000000000000000000000000, `__LINE__); //   8: fn=SHR, a=0X00000000, b= 2, y=0X00000000
	test_case({2'b11, 32'b00000000000000000000000000000000, 5'b00010}, 32'b00000000000000000000000000000000, `__LINE__); //   9: fn=SRA, a=0X00000000, b= 2, y=0X00000000
	test_case({2'b00, 32'b00000000000000000000000000000000, 5'b00100}, 32'b00000000000000000000000000000000, `__LINE__); //  10: fn=SHL, a=0X00000000, b= 4, y=0X00000000
	test_case({2'b01, 32'b00000000000000000000000000000000, 5'b00100}, 32'b00000000000000000000000000000000, `__LINE__); //  11: fn=SHR, a=0X00000000, b= 4, y=0X00000000
	test_case({2'b11, 32'b00000000000000000000000000000000, 5'b00100}, 32'b00000000000000000000000000000000, `__LINE__); //  12: fn=SRA, a=0X00000000, b= 4, y=0X00000000
	test_case({2'b00, 32'b00000000000000000000000000000000, 5'b01000}, 32'b00000000000000000000000000000000, `__LINE__); //  13: fn=SHL, a=0X00000000, b= 8, y=0X00000000
	test_case({2'b01, 32'b00000000000000000000000000000000, 5'b01000}, 32'b00000000000000000000000000000000, `__LINE__); //  14: fn=SHR, a=0X00000000, b= 8, y=0X00000000
	test_case({2'b11, 32'b00000000000000000000000000000000, 5'b01000}, 32'b00000000000000000000000000000000, `__LINE__); //  15: fn=SRA, a=0X00000000, b= 8, y=0X00000000
	test_case({2'b00, 32'b00000000000000000000000000000000, 5'b10000}, 32'b00000000000000000000000000000000, `__LINE__); //  16: fn=SHL, a=0X00000000, b=16, y=0X00000000
	test_case({2'b01, 32'b00000000000000000000000000000000, 5'b10000}, 32'b00000000000000000000000000000000, `__LINE__); //  17: fn=SHR, a=0X00000000, b=16, y=0X00000000
	test_case({2'b11, 32'b00000000000000000000000000000000, 5'b10000}, 32'b00000000000000000000000000000000, `__LINE__); //  18: fn=SRA, a=0X00000000, b=16, y=0X00000000
	test_case({2'b00, 32'b00000000000000000000000000000000, 5'b11111}, 32'b00000000000000000000000000000000, `__LINE__); //  19: fn=SHL, a=0X00000000, b=31, y=0X00000000
	test_case({2'b01, 32'b00000000000000000000000000000000, 5'b11111}, 32'b00000000000000000000000000000000, `__LINE__); //  20: fn=SHR, a=0X00000000, b=31, y=0X00000000
	test_case({2'b11, 32'b00000000000000000000000000000000, 5'b11111}, 32'b00000000000000000000000000000000, `__LINE__); //  21: fn=SRA, a=0X00000000, b=31, y=0X00000000
	test_case({2'b00, 32'b00000000000000000000000000000001, 5'b00000}, 32'b00000000000000000000000000000001, `__LINE__); //  22: fn=SHL, a=0X00000001, b= 0, y=0X00000001
	test_case({2'b01, 32'b00000000000000000000000000000001, 5'b00000}, 32'b00000000000000000000000000000001, `__LINE__); //  23: fn=SHR, a=0X00000001, b= 0, y=0X00000001
	test_case({2'b11, 32'b00000000000000000000000000000001, 5'b00000}, 32'b00000000000000000000000000000001, `__LINE__); //  24: fn=SRA, a=0X00000001, b= 0, y=0X00000001
	test_case({2'b00, 32'b00000000000000000000000000000001, 5'b00001}, 32'b00000000000000000000000000000010, `__LINE__); //  25: fn=SHL, a=0X00000001, b= 1, y=0X00000002
	test_case({2'b01, 32'b00000000000000000000000000000001, 5'b00001}, 32'b00000000000000000000000000000000, `__LINE__); //  26: fn=SHR, a=0X00000001, b= 1, y=0X00000000
	test_case({2'b11, 32'b00000000000000000000000000000001, 5'b00001}, 32'b00000000000000000000000000000000, `__LINE__); //  27: fn=SRA, a=0X00000001, b= 1, y=0X00000000
	test_case({2'b00, 32'b00000000000000000000000000000001, 5'b00010}, 32'b00000000000000000000000000000100, `__LINE__); //  28: fn=SHL, a=0X00000001, b= 2, y=0X00000004
	test_case({2'b01, 32'b00000000000000000000000000000001, 5'b00010}, 32'b00000000000000000000000000000000, `__LINE__); //  29: fn=SHR, a=0X00000001, b= 2, y=0X00000000
	test_case({2'b11, 32'b00000000000000000000000000000001, 5'b00010}, 32'b00000000000000000000000000000000, `__LINE__); //  30: fn=SRA, a=0X00000001, b= 2, y=0X00000000
	test_case({2'b00, 32'b00000000000000000000000000000001, 5'b00100}, 32'b00000000000000000000000000010000, `__LINE__); //  31: fn=SHL, a=0X00000001, b= 4, y=0X00000010
	test_case({2'b01, 32'b00000000000000000000000000000001, 5'b00100}, 32'b00000000000000000000000000000000, `__LINE__); //  32: fn=SHR, a=0X00000001, b= 4, y=0X00000000
	test_case({2'b11, 32'b00000000000000000000000000000001, 5'b00100}, 32'b00000000000000000000000000000000, `__LINE__); //  33: fn=SRA, a=0X00000001, b= 4, y=0X00000000
	test_case({2'b00, 32'b00000000000000000000000000000001, 5'b01000}, 32'b00000000000000000000000100000000, `__LINE__); //  34: fn=SHL, a=0X00000001, b= 8, y=0X00000100
	test_case({2'b01, 32'b00000000000000000000000000000001, 5'b01000}, 32'b00000000000000000000000000000000, `__LINE__); //  35: fn=SHR, a=0X00000001, b= 8, y=0X00000000
	test_case({2'b11, 32'b00000000000000000000000000000001, 5'b01000}, 32'b00000000000000000000000000000000, `__LINE__); //  36: fn=SRA, a=0X00000001, b= 8, y=0X00000000
	test_case({2'b00, 32'b00000000000000000000000000000001, 5'b10000}, 32'b00000000000000010000000000000000, `__LINE__); //  37: fn=SHL, a=0X00000001, b=16, y=0X00010000
	test_case({2'b01, 32'b00000000000000000000000000000001, 5'b10000}, 32'b00000000000000000000000000000000, `__LINE__); //  38: fn=SHR, a=0X00000001, b=16, y=0X00000000
	test_case({2'b11, 32'b00000000000000000000000000000001, 5'b10000}, 32'b00000000000000000000000000000000, `__LINE__); //  39: fn=SRA, a=0X00000001, b=16, y=0X00000000
	test_case({2'b00, 32'b00000000000000000000000000000001, 5'b11111}, 32'b10000000000000000000000000000000, `__LINE__); //  40: fn=SHL, a=0X00000001, b=31, y=0X80000000
	test_case({2'b01, 32'b00000000000000000000000000000001, 5'b11111}, 32'b00000000000000000000000000000000, `__LINE__); //  41: fn=SHR, a=0X00000001, b=31, y=0X00000000
	test_case({2'b11, 32'b00000000000000000000000000000001, 5'b11111}, 32'b00000000000000000000000000000000, `__LINE__); //  42: fn=SRA, a=0X00000001, b=31, y=0X00000000
	test_case({2'b00, 32'b11111111111111111111111111111111, 5'b00000}, 32'b11111111111111111111111111111111, `__LINE__); //  43: fn=SHL, a=0XFFFFFFFF, b= 0, y=0XFFFFFFFF
	test_case({2'b01, 32'b11111111111111111111111111111111, 5'b00000}, 32'b11111111111111111111111111111111, `__LINE__); //  44: fn=SHR, a=0XFFFFFFFF, b= 0, y=0XFFFFFFFF
	test_case({2'b11, 32'b11111111111111111111111111111111, 5'b00000}, 32'b11111111111111111111111111111111, `__LINE__); //  45: fn=SRA, a=0XFFFFFFFF, b= 0, y=0XFFFFFFFF
	test_case({2'b00, 32'b11111111111111111111111111111111, 5'b00001}, 32'b11111111111111111111111111111110, `__LINE__); //  46: fn=SHL, a=0XFFFFFFFF, b= 1, y=0XFFFFFFFE
	test_case({2'b01, 32'b11111111111111111111111111111111, 5'b00001}, 32'b01111111111111111111111111111111, `__LINE__); //  47: fn=SHR, a=0XFFFFFFFF, b= 1, y=0X7FFFFFFF
	test_case({2'b11, 32'b11111111111111111111111111111111, 5'b00001}, 32'b11111111111111111111111111111111, `__LINE__); //  48: fn=SRA, a=0XFFFFFFFF, b= 1, y=0XFFFFFFFF
	test_case({2'b00, 32'b11111111111111111111111111111111, 5'b00010}, 32'b11111111111111111111111111111100, `__LINE__); //  49: fn=SHL, a=0XFFFFFFFF, b= 2, y=0XFFFFFFFC
	test_case({2'b01, 32'b11111111111111111111111111111111, 5'b00010}, 32'b00111111111111111111111111111111, `__LINE__); //  50: fn=SHR, a=0XFFFFFFFF, b= 2, y=0X3FFFFFFF
	test_case({2'b11, 32'b11111111111111111111111111111111, 5'b00010}, 32'b11111111111111111111111111111111, `__LINE__); //  51: fn=SRA, a=0XFFFFFFFF, b= 2, y=0XFFFFFFFF
	test_case({2'b00, 32'b11111111111111111111111111111111, 5'b00100}, 32'b11111111111111111111111111110000, `__LINE__); //  52: fn=SHL, a=0XFFFFFFFF, b= 4, y=0XFFFFFFF0
	test_case({2'b01, 32'b11111111111111111111111111111111, 5'b00100}, 32'b00001111111111111111111111111111, `__LINE__); //  53: fn=SHR, a=0XFFFFFFFF, b= 4, y=0X0FFFFFFF
	test_case({2'b11, 32'b11111111111111111111111111111111, 5'b00100}, 32'b11111111111111111111111111111111, `__LINE__); //  54: fn=SRA, a=0XFFFFFFFF, b= 4, y=0XFFFFFFFF
	test_case({2'b00, 32'b11111111111111111111111111111111, 5'b01000}, 32'b11111111111111111111111100000000, `__LINE__); //  55: fn=SHL, a=0XFFFFFFFF, b= 8, y=0XFFFFFF00
	test_case({2'b01, 32'b11111111111111111111111111111111, 5'b01000}, 32'b00000000111111111111111111111111, `__LINE__); //  56: fn=SHR, a=0XFFFFFFFF, b= 8, y=0X00FFFFFF
	test_case({2'b11, 32'b11111111111111111111111111111111, 5'b01000}, 32'b11111111111111111111111111111111, `__LINE__); //  57: fn=SRA, a=0XFFFFFFFF, b= 8, y=0XFFFFFFFF
	test_case({2'b00, 32'b11111111111111111111111111111111, 5'b10000}, 32'b11111111111111110000000000000000, `__LINE__); //  58: fn=SHL, a=0XFFFFFFFF, b=16, y=0XFFFF0000
	test_case({2'b01, 32'b11111111111111111111111111111111, 5'b10000}, 32'b00000000000000001111111111111111, `__LINE__); //  59: fn=SHR, a=0XFFFFFFFF, b=16, y=0X0000FFFF
	test_case({2'b11, 32'b11111111111111111111111111111111, 5'b10000}, 32'b11111111111111111111111111111111, `__LINE__); //  60: fn=SRA, a=0XFFFFFFFF, b=16, y=0XFFFFFFFF
	test_case({2'b00, 32'b11111111111111111111111111111111, 5'b11111}, 32'b10000000000000000000000000000000, `__LINE__); //  61: fn=SHL, a=0XFFFFFFFF, b=31, y=0X80000000
	test_case({2'b01, 32'b11111111111111111111111111111111, 5'b11111}, 32'b00000000000000000000000000000001, `__LINE__); //  62: fn=SHR, a=0XFFFFFFFF, b=31, y=0X00000001
	test_case({2'b11, 32'b11111111111111111111111111111111, 5'b11111}, 32'b11111111111111111111111111111111, `__LINE__); //  63: fn=SRA, a=0XFFFFFFFF, b=31, y=0XFFFFFFFF
	test_case({2'b00, 32'b00010010001101000101011001111000, 5'b00000}, 32'b00010010001101000101011001111000, `__LINE__); //  64: fn=SHL, a=0X12345678, b= 0, y=0X12345678
	test_case({2'b01, 32'b00010010001101000101011001111000, 5'b00000}, 32'b00010010001101000101011001111000, `__LINE__); //  65: fn=SHR, a=0X12345678, b= 0, y=0X12345678
	test_case({2'b11, 32'b00010010001101000101011001111000, 5'b00000}, 32'b00010010001101000101011001111000, `__LINE__); //  66: fn=SRA, a=0X12345678, b= 0, y=0X12345678
	test_case({2'b00, 32'b00010010001101000101011001111000, 5'b00001}, 32'b00100100011010001010110011110000, `__LINE__); //  67: fn=SHL, a=0X12345678, b= 1, y=0X2468ACF0
	test_case({2'b01, 32'b00010010001101000101011001111000, 5'b00001}, 32'b00001001000110100010101100111100, `__LINE__); //  68: fn=SHR, a=0X12345678, b= 1, y=0X091A2B3C
	test_case({2'b11, 32'b00010010001101000101011001111000, 5'b00001}, 32'b00001001000110100010101100111100, `__LINE__); //  69: fn=SRA, a=0X12345678, b= 1, y=0X091A2B3C
	test_case({2'b00, 32'b00010010001101000101011001111000, 5'b00010}, 32'b01001000110100010101100111100000, `__LINE__); //  70: fn=SHL, a=0X12345678, b= 2, y=0X48D159E0
	test_case({2'b01, 32'b00010010001101000101011001111000, 5'b00010}, 32'b00000100100011010001010110011110, `__LINE__); //  71: fn=SHR, a=0X12345678, b= 2, y=0X048D159E
	test_case({2'b11, 32'b00010010001101000101011001111000, 5'b00010}, 32'b00000100100011010001010110011110, `__LINE__); //  72: fn=SRA, a=0X12345678, b= 2, y=0X048D159E
	test_case({2'b00, 32'b00010010001101000101011001111000, 5'b00100}, 32'b00100011010001010110011110000000, `__LINE__); //  73: fn=SHL, a=0X12345678, b= 4, y=0X23456780
	test_case({2'b01, 32'b00010010001101000101011001111000, 5'b00100}, 32'b00000001001000110100010101100111, `__LINE__); //  74: fn=SHR, a=0X12345678, b= 4, y=0X01234567
	test_case({2'b11, 32'b00010010001101000101011001111000, 5'b00100}, 32'b00000001001000110100010101100111, `__LINE__); //  75: fn=SRA, a=0X12345678, b= 4, y=0X01234567
	test_case({2'b00, 32'b00010010001101000101011001111000, 5'b01000}, 32'b00110100010101100111100000000000, `__LINE__); //  76: fn=SHL, a=0X12345678, b= 8, y=0X34567800
	test_case({2'b01, 32'b00010010001101000101011001111000, 5'b01000}, 32'b00000000000100100011010001010110, `__LINE__); //  77: fn=SHR, a=0X12345678, b= 8, y=0X00123456
	test_case({2'b11, 32'b00010010001101000101011001111000, 5'b01000}, 32'b00000000000100100011010001010110, `__LINE__); //  78: fn=SRA, a=0X12345678, b= 8, y=0X00123456
	test_case({2'b00, 32'b00010010001101000101011001111000, 5'b10000}, 32'b01010110011110000000000000000000, `__LINE__); //  79: fn=SHL, a=0X12345678, b=16, y=0X56780000
	test_case({2'b01, 32'b00010010001101000101011001111000, 5'b10000}, 32'b00000000000000000001001000110100, `__LINE__); //  80: fn=SHR, a=0X12345678, b=16, y=0X00001234
	test_case({2'b11, 32'b00010010001101000101011001111000, 5'b10000}, 32'b00000000000000000001001000110100, `__LINE__); //  81: fn=SRA, a=0X12345678, b=16, y=0X00001234
	test_case({2'b00, 32'b00010010001101000101011001111000, 5'b11111}, 32'b00000000000000000000000000000000, `__LINE__); //  82: fn=SHL, a=0X12345678, b=31, y=0X00000000
	test_case({2'b01, 32'b00010010001101000101011001111000, 5'b11111}, 32'b00000000000000000000000000000000, `__LINE__); //  83: fn=SHR, a=0X12345678, b=31, y=0X00000000
	test_case({2'b11, 32'b00010010001101000101011001111000, 5'b11111}, 32'b00000000000000000000000000000000, `__LINE__); //  84: fn=SRA, a=0X12345678, b=31, y=0X00000000
	test_case({2'b00, 32'b11111110110111001011101010011000, 5'b00000}, 32'b11111110110111001011101010011000, `__LINE__); //  85: fn=SHL, a=0XFEDCBA98, b= 0, y=0XFEDCBA98
	test_case({2'b01, 32'b11111110110111001011101010011000, 5'b00000}, 32'b11111110110111001011101010011000, `__LINE__); //  86: fn=SHR, a=0XFEDCBA98, b= 0, y=0XFEDCBA98
	test_case({2'b11, 32'b11111110110111001011101010011000, 5'b00000}, 32'b11111110110111001011101010011000, `__LINE__); //  87: fn=SRA, a=0XFEDCBA98, b= 0, y=0XFEDCBA98
	test_case({2'b00, 32'b11111110110111001011101010011000, 5'b00001}, 32'b11111101101110010111010100110000, `__LINE__); //  88: fn=SHL, a=0XFEDCBA98, b= 1, y=0XFDB97530
	test_case({2'b01, 32'b11111110110111001011101010011000, 5'b00001}, 32'b01111111011011100101110101001100, `__LINE__); //  89: fn=SHR, a=0XFEDCBA98, b= 1, y=0X7F6E5D4C
	test_case({2'b11, 32'b11111110110111001011101010011000, 5'b00001}, 32'b11111111011011100101110101001100, `__LINE__); //  90: fn=SRA, a=0XFEDCBA98, b= 1, y=0XFF6E5D4C
	test_case({2'b00, 32'b11111110110111001011101010011000, 5'b00010}, 32'b11111011011100101110101001100000, `__LINE__); //  91: fn=SHL, a=0XFEDCBA98, b= 2, y=0XFB72EA60
	test_case({2'b01, 32'b11111110110111001011101010011000, 5'b00010}, 32'b00111111101101110010111010100110, `__LINE__); //  92: fn=SHR, a=0XFEDCBA98, b= 2, y=0X3FB72EA6
	test_case({2'b11, 32'b11111110110111001011101010011000, 5'b00010}, 32'b11111111101101110010111010100110, `__LINE__); //  93: fn=SRA, a=0XFEDCBA98, b= 2, y=0XFFB72EA6
	test_case({2'b00, 32'b11111110110111001011101010011000, 5'b00100}, 32'b11101101110010111010100110000000, `__LINE__); //  94: fn=SHL, a=0XFEDCBA98, b= 4, y=0XEDCBA980
	test_case({2'b01, 32'b11111110110111001011101010011000, 5'b00100}, 32'b00001111111011011100101110101001, `__LINE__); //  95: fn=SHR, a=0XFEDCBA98, b= 4, y=0X0FEDCBA9
	test_case({2'b11, 32'b11111110110111001011101010011000, 5'b00100}, 32'b11111111111011011100101110101001, `__LINE__); //  96: fn=SRA, a=0XFEDCBA98, b= 4, y=0XFFEDCBA9
	test_case({2'b00, 32'b11111110110111001011101010011000, 5'b01000}, 32'b11011100101110101001100000000000, `__LINE__); //  97: fn=SHL, a=0XFEDCBA98, b= 8, y=0XDCBA9800
	test_case({2'b01, 32'b11111110110111001011101010011000, 5'b01000}, 32'b00000000111111101101110010111010, `__LINE__); //  98: fn=SHR, a=0XFEDCBA98, b= 8, y=0X00FEDCBA
	test_case({2'b11, 32'b11111110110111001011101010011000, 5'b01000}, 32'b11111111111111101101110010111010, `__LINE__); //  99: fn=SRA, a=0XFEDCBA98, b= 8, y=0XFFFEDCBA
	test_case({2'b00, 32'b11111110110111001011101010011000, 5'b10000}, 32'b10111010100110000000000000000000, `__LINE__); // 100: fn=SHL, a=0XFEDCBA98, b=16, y=0XBA980000
	test_case({2'b01, 32'b11111110110111001011101010011000, 5'b10000}, 32'b00000000000000001111111011011100, `__LINE__); // 101: fn=SHR, a=0XFEDCBA98, b=16, y=0X0000FEDC
	test_case({2'b11, 32'b11111110110111001011101010011000, 5'b10000}, 32'b11111111111111111111111011011100, `__LINE__); // 102: fn=SRA, a=0XFEDCBA98, b=16, y=0XFFFFFEDC
	test_case({2'b00, 32'b11111110110111001011101010011000, 5'b11111}, 32'b00000000000000000000000000000000, `__LINE__); // 103: fn=SHL, a=0XFEDCBA98, b=31, y=0X00000000
	test_case({2'b01, 32'b11111110110111001011101010011000, 5'b11111}, 32'b00000000000000000000000000000001, `__LINE__); // 104: fn=SHR, a=0XFEDCBA98, b=31, y=0X00000001
	test_case({2'b11, 32'b11111110110111001011101010011000, 5'b11111}, 32'b11111111111111111111111111111111, `__LINE__); // 105: fn=SRA, a=0XFEDCBA98, b=31, y=0XFFFFFFFF
	$display("");
	if (dut_error != 0) begin
		$display("ERROR: %d test cases failed", dut_error);
		$finish_and_return(1);
	end
	$display("PASS:  all test cases passed");
	$display("");
    $finish;
end


alu_shift dut (
    .sfn(sfn),
    .a(a),
    .b(b),
    .y(y)
);

endmodule
