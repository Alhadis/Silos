module design(I1,I2,I3,I4,I5,I6,I7,I8,I9,I10,I11,I12,I13,I14,I15,I16,I17,I18,I19,I20,I21,I22,I23,I24,I25,I26,I27,I28,I29,O1,O2,O3,O4,O5,O6,O7);
input I1;
input I2;
input I3;
input I4;
input I5;
input I6;
input I7;
input I8;
input I9;
input I10;
input I11;
input I12;
input I13;
input I14;
input I15;
input I16;
input I17;
input I18;
input I19;
input I20;
input I21;
input I22;
input I23;
input I24;
input I25;
input I26;
input I27;
input I28;
input I29;

output O1;
output O2;
output O3;
output O4;
output O5;
output O6;
output O7;

wire W1;
wire W2;
wire W3;
wire W4;
wire W5;
wire W6;
wire W7;
wire W8;
wire W9;
wire W10;
wire W11;
wire W12;
wire W13;
wire W14;
wire W15;
wire W16;
wire W17;
wire W18;
wire W19;
wire W20;
wire W21;
wire W22;
wire W23;
wire W24;
wire W25;
wire W26;
wire W27;
wire W28;
wire W29;
wire W30;
wire W31;
wire W32;
wire W33;
wire W34;
wire W35;
wire W36;
wire W37;
wire W38;
wire W39;
wire W40;
wire W41;
wire W42;
wire W43;
wire W44;
wire W45;
wire W46;
wire W47;
wire W48;
wire W49;
wire W50;
wire W51;
wire W52;
wire W53;
wire W54;
wire W55;
wire W56;
wire W57;
wire W58;
wire W59;
wire W60;
wire W61;
wire W62;
wire W63;
wire W64;
wire W65;
wire W66;
wire W67;
wire W68;
wire W69;
wire W70;
wire W71;
wire W72;
wire W73;
wire W74;
wire W75;
wire W76;
wire W77;
wire W78;
wire W79;
wire W80;
wire W81;
wire W82;
wire W83;
wire W84;
wire W85;
wire W86;
wire W87;
wire W88;
wire W89;
wire W90;
wire W91;
wire W92;
wire W93;
wire W94;
wire W95;
wire W96;
wire W97;
wire W98;
wire W99;
wire W100;
wire W101;
wire W102;
wire W103;
wire W104;
wire W105;
wire W106;
wire W107;
wire W108;
wire W109;
wire W110;
wire W111;
wire W112;
wire W113;
wire W114;
wire W115;
wire W116;
wire W117;
wire W118;
wire W119;
wire W120;
wire W121;
wire W122;
wire W123;
wire W124;
wire W125;
wire W126;
wire W127;
wire W128;
wire W129;
wire W130;
wire W131;
wire W132;
wire W133;
wire W134;
wire W135;
wire W136;
wire W137;
wire W138;
wire W139;
wire W140;
wire W141;
wire W142;
wire W143;
wire W144;
wire W145;
wire W146;
wire W147;
wire W148;
wire W149;
wire W150;
wire W151;
wire W152;
wire W153;
wire W154;
wire W155;
wire W156;
wire W157;
wire W158;
wire W159;
wire W160;
wire W161;
wire W162;
wire W163;
wire W164;
wire W165;
wire W166;
wire W167;
wire W168;
wire W169;
wire W170;
wire W171;
wire W172;
wire W173;
wire W174;
wire W175;
wire W176;
wire W177;
wire W178;
wire W179;
wire W180;
wire W181;
wire W182;
wire W183;
wire W184;
wire W185;
wire W186;
wire W187;
wire W188;
wire W189;
wire W190;
wire W191;
wire W192;
wire W193;
wire W194;
wire W195;
wire W196;
wire W197;
wire W198;
wire W199;
wire W200;
wire W201;
wire W202;
wire W203;
wire W204;
wire W205;
wire W206;
wire W207;
wire W208;
wire W209;
wire W210;
wire W211;
wire W212;
wire W213;
wire W214;
wire W215;
wire W216;
wire W217;
wire W218;
wire W219;
wire W220;
wire W221;
wire W222;
wire W223;
wire W224;
wire W225;
wire W226;
wire W227;
wire W228;
wire W229;
wire W230;
wire W231;
wire W232;
wire W233;
wire W234;
wire W235;
wire W236;
wire W237;
wire W238;
wire W239;
wire W240;
wire W241;
wire W242;
wire W243;
wire W244;
wire W245;
wire W246;
wire W247;
wire W248;
wire W249;
wire W250;
wire W251;
wire W252;
wire W253;
wire W254;
wire W255;
wire W256;
wire W257;
wire W258;
wire W259;
wire W260;
wire W261;
wire W262;
wire W263;
wire W264;
wire W265;
wire W266;
wire W267;
wire W268;
wire W269;
wire W270;
wire W271;
wire W272;
wire W273;
wire W274;
wire W275;
wire W276;
wire W277;
wire W278;
wire W279;
wire W280;
wire W281;
wire W282;
wire W283;
wire W284;
wire W285;
wire W286;
wire W287;
wire W288;
wire W289;
wire W290;
wire W291;
wire W292;
wire W293;
wire W294;
wire W295;
wire W296;
wire W297;
wire W298;
wire W299;
wire W300;
wire W301;
wire W302;
wire W303;
wire W304;
wire W305;
wire W306;
wire W307;
wire W308;
wire W309;
wire W310;
wire W311;
wire W312;
wire W313;
wire W314;
wire W315;
wire W316;
wire W317;
wire W318;
wire W319;
wire W320;
wire W321;
wire W322;
wire W323;
wire W324;
wire W325;
wire W326;
wire W327;
wire W328;
wire W329;
wire W330;
wire W331;
wire W332;
wire W333;
wire W334;
wire W335;
wire W336;
wire W337;
wire W338;
wire W339;
wire W340;
wire W341;
wire W342;
wire W343;
wire W344;
wire W345;
wire W346;
wire W347;
wire W348;
wire W349;
wire W350;
wire W351;

not G1 (O1, W1);
not G2 (O2, W2);
not G3 (O3, W3);
not G4 (O4, W4);
not G5 (O5, W5);
not G6 (O6, W6);
not G7 (O7, W7);
not G8 (W1, W8);
not G9 (W2, W9);
not G10 (W3, W10);
not G11 (W4, W11);
not G12 (W5, W12);
not G13 (W6, W13);
not G14 (W7, W14);
not G15 (W8, W15);
not G16 (W9, W16);
not G17 (W10, W17);
not G18 (W11, W18);
not G19 (W12, W19);
not G20 (W13, W20);
not G21 (W14, W21);
not G22 (W15, W22);
not G23 (W16, W23);
not G24 (W17, W24);
not G25 (W18, W25);
not G26 (W19, W26);
not G27 (W20, W27);
not G28 (W21, W28);
or G29 (W22, W29, W30);
or G30 (W23, W31, W32);
or G31 (W24, W33, W34);
or G32 (W25, W35, W36);
or G33 (W26, W37, W38);
or G34 (W27, W39, W40);
or G35 (W28, W41, W42);
and G36 (W29, W43, W44);
and G37 (W30, W45, W46);
and G38 (W31, W47, W48);
and G39 (W32, W49, W50);
and G40 (W33, W51, W52);
and G41 (W34, W53, W54);
and G42 (W35, W55, W56);
and G43 (W36, W57, W58);
and G44 (W37, W59, W60);
and G45 (W38, W61, W62);
and G46 (W39, W63, W64);
and G47 (W40, W65, W66);
and G48 (W41, W67, W68);
and G49 (W42, W69, W70);
or G50 (W43, W71, W72);
not G51 (W44, W46);
not G52 (W45, W73);
not G53 (W46, W74);
or G54 (W47, W75, W76);
not G55 (W48, W50);
not G56 (W49, W77);
not G57 (W50, W78);
or G58 (W51, W79, W80);
not G59 (W52, W54);
not G60 (W53, W81);
not G61 (W54, W82);
or G62 (W55, W83, W84);
not G63 (W56, W58);
not G64 (W57, W85);
not G65 (W58, W86);
or G66 (W59, W87, W88);
not G67 (W60, W62);
not G68 (W61, W89);
not G69 (W62, W90);
or G70 (W63, W91, W92);
not G71 (W64, W66);
not G72 (W65, W93);
not G73 (W66, W94);
or G74 (W67, W95, W96);
not G75 (W68, W70);
not G76 (W69, W97);
not G77 (W70, W98);
and G78 (W71, I1, W99);
and G79 (W72, W100, W101);
not G80 (W73, W102);
not G81 (W74, W103);
and G82 (W75, I2, W104);
and G83 (W76, W105, W106);
not G84 (W77, W107);
not G85 (W78, W103);
and G86 (W79, I3, W108);
and G87 (W80, W109, W110);
not G88 (W81, W111);
not G89 (W82, W103);
and G90 (W83, I4, W112);
and G91 (W84, W113, W114);
not G92 (W85, W115);
not G93 (W86, W103);
and G94 (W87, I5, W116);
and G95 (W88, W117, W118);
not G96 (W89, W119);
not G97 (W90, W103);
and G98 (W91, I6, W120);
and G99 (W92, W121, W122);
not G100 (W93, W123);
not G101 (W94, W103);
and G102 (W95, I7, W124);
and G103 (W96, W125, W126);
not G104 (W97, W127);
not G105 (W98, W103);
not G106 (W99, W101);
nand G107 (W100, W128, W129);
not G108 (W101, W130);
not G109 (W102, W131);
or G110 (W103, W132, W133);
not G111 (W104, W106);
nand G112 (W105, W134, W135);
not G113 (W106, W136);
not G114 (W107, W137);
not G115 (W108, W110);
nand G116 (W109, W138, W139);
not G117 (W110, W140);
not G118 (W111, W141);
not G119 (W112, W114);
nand G120 (W113, W142, W143);
not G121 (W114, W144);
not G122 (W115, W145);
not G123 (W116, W118);
nand G124 (W117, W146, W147);
not G125 (W118, W148);
not G126 (W119, W149);
not G127 (W120, W122);
nand G128 (W121, W150, W151);
not G129 (W122, W152);
not G130 (W123, W153);
not G131 (W124, W126);
nand G132 (W125, W154, W155);
not G133 (W126, W156);
not G134 (W127, W157);
nand G135 (W128, I1, W158);
nand G136 (W129, W159, W158);
not G137 (W130, W160);
not G138 (W131, W161);
not G139 (W132, W162);
and G140 (W133, W163, W164);
nand G141 (W134, I2, W165);
nand G142 (W135, W166, W165);
not G143 (W136, W160);
not G144 (W137, W167);
nand G145 (W138, I3, W168);
nand G146 (W139, W169, W168);
not G147 (W140, W160);
not G148 (W141, W170);
nand G149 (W142, I4, W171);
nand G150 (W143, W172, W171);
not G151 (W144, W160);
not G152 (W145, W173);
nand G153 (W146, I5, W174);
nand G154 (W147, W175, W174);
not G155 (W148, W160);
not G156 (W149, W176);
nand G157 (W150, I6, W177);
nand G158 (W151, W178, W177);
not G159 (W152, W160);
not G160 (W153, W179);
nand G161 (W154, I7, W180);
nand G162 (W155, W181, W180);
not G163 (W156, W160);
not G164 (W157, W182);
nand G165 (W158, I1, W159);
or G166 (W159, W183, W184);
or G167 (W160, W164, W185);
not G168 (W161, W186);
not G169 (W162, W187);
or G170 (W163, W188, W189);
or G171 (W164, W190, W191);
nand G172 (W165, I2, W166);
or G173 (W166, W192, W193);
not G174 (W167, W194);
nand G175 (W168, I3, W169);
or G176 (W169, W195, W196);
not G177 (W170, W197);
nand G178 (W171, I4, W172);
or G179 (W172, W198, W199);
not G180 (W173, W200);
nand G181 (W174, I5, W175);
or G182 (W175, W201, W202);
not G183 (W176, W203);
nand G184 (W177, I6, W178);
or G185 (W178, W204, W205);
not G186 (W179, W206);
nand G187 (W180, I7, W181);
or G188 (W181, W207, W208);
not G189 (W182, W209);
and G190 (W183, W210, W211);
and G191 (W184, I8, W212);
not G192 (W185, W213);
not G193 (W186, W214);
not G194 (W187, W215);
and G195 (W188, W216, W217);
and G196 (W189, W218, W219);
and G197 (W190, W220, W221);
and G198 (W191, W222, W223);
and G199 (W192, W224, W225);
and G200 (W193, I9, W226);
not G201 (W194, W227);
and G202 (W195, W228, W229);
and G203 (W196, I10, W230);
not G204 (W197, W231);
not G205 (W198, W232);
and G206 (W199, I11, W233);
not G207 (W200, W234);
and G208 (W201, W235, W236);
and G209 (W202, I12, W237);
not G210 (W203, W238);
and G211 (W204, W239, W240);
and G212 (W205, I13, W241);
not G213 (W206, W242);
and G214 (W207, W243, W244);
and G215 (W208, I14, W245);
not G216 (W209, W246);
or G217 (W210, W247, W248);
not G218 (W211, W212);
not G219 (W212, W249);
not G220 (W213, W250);
not G221 (W214, W251);
nand G222 (W215, W252, W253, W254);
and G223 (W216, W255, W256);
not G224 (W217, W219);
and G225 (W218, W257, I6);
not G226 (W219, W258);
nand G227 (W220, W253, W259);
and G228 (W221, W223, I15);
not G229 (W222, W260);
and G230 (W223, W261, W262);
or G231 (W224, W263, W264);
not G232 (W225, W226);
not G233 (W226, W265);
not G234 (W227, W251);
or G235 (W228, W266, W267);
not G236 (W229, W230);
not G237 (W230, W268);
not G238 (W231, W251);
not G239 (W232, W269);
not G240 (W233, W270);
not G241 (W234, W251);
or G242 (W235, W271, W272);
not G243 (W236, W237);
not G244 (W237, W273);
not G245 (W238, W251);
or G246 (W239, W274, W275);
not G247 (W240, W241);
not G248 (W241, W276);
not G249 (W242, W251);
or G250 (W243, W277, W278);
not G251 (W244, W245);
not G252 (W245, W279);
not G253 (W246, W251);
and G254 (W247, W280, W281);
and G255 (W248, W282, W283);
not G256 (W249, W185);
nand G257 (W250, W284, W285);
or G258 (W251, W286, W132);
not G259 (W252, I16);
not G260 (W253, I17);
and G261 (W254, W287, W259);
and G262 (W255, W288, W289);
not G263 (W256, I6);
and G264 (W257, W290, I3);
not G265 (W258, W291);
not G266 (W259, I18);
nand G267 (W260, W292, I16, I19);
not G268 (W261, W293);
and G269 (W262, W294, W295);
and G270 (W263, W296, W297);
and G271 (W264, W298, W299);
not G272 (W265, W185);
and G273 (W266, W288, W300);
and G274 (W267, W290, W301);
not G275 (W268, W185);
not G276 (W269, W233);
not G277 (W270, W185);
and G278 (W271, W302, W303);
and G279 (W272, W304, W305);
not G280 (W273, W185);
and G281 (W274, W255, W306);
and G282 (W275, W257, W307);
not G283 (W276, W185);
and G284 (W277, W308, W309);
and G285 (W278, W310, W311);
not G286 (W279, W185);
and G287 (W280, W312, W313);
not G288 (W281, W283);
and G289 (W282, W314, I20);
not G290 (W283, W315);
nand G291 (W284, W316, W223);
nand G292 (W285, I21, W223);
nand G293 (W286, W317, W318);
not G294 (W287, I19);
and G295 (W288, W319, W320);
not G296 (W289, I3);
and G297 (W290, W321, I22);
not G298 (W291, W322);
not G299 (W292, I21);
not G300 (W293, W323);
not G301 (W294, I23);
and G302 (W295, W324, W325);
and G303 (W296, W280, W326);
not G304 (W297, W299);
and G305 (W298, W282, I1);
not G306 (W299, W327);
not G307 (W300, W301);
not G308 (W301, W328);
and G309 (W302, W308, W329);
not G310 (W303, W305);
and G311 (W304, W310, I7);
not G312 (W305, W330);
not G313 (W306, W307);
not G314 (W307, W331);
not G315 (W308, W332);
not G316 (W309, W311);
not G317 (W310, W333);
not G318 (W311, W334);
and G319 (W312, W302, W335);
not G320 (W313, I20);
and G321 (W314, W304, I5);
not G322 (W315, W291);
not G323 (W316, W336);
and G324 (W317, W337, W260);
nand G325 (W318, I18, W252, W253);
and G326 (W319, W296, W338);
not G327 (W320, I22);
and G328 (W321, W298, I2);
not G329 (W322, W339);
not G330 (W323, W340);
not G331 (W324, I24);
and G332 (W325, W341, W342);
not G333 (W326, I1);
not G334 (W327, W291);
not G335 (W328, W291);
not G336 (W329, I7);
not G337 (W330, W291);
not G338 (W331, W291);
not G339 (W332, W343);
not G340 (W333, I4);
not G341 (W334, W291);
not G342 (W335, I5);
nand G343 (W336, W344, W292, W254);
nand G344 (W337, I17, W259);
not G345 (W338, I2);
nand G346 (W339, W345, W318, W346);
not G347 (W340, I25);
not G348 (W341, I26);
and G349 (W342, W347, W348);
not G350 (W343, I4);
not G351 (W344, W345);
nand G352 (W345, I16, W253);
nand G353 (W346, W349, W252);
not G354 (W347, I27);
and G355 (W348, W350, W351);
not G356 (W349, W337);
not G357 (W350, I28);
not G358 (W351, I29);
endmodule