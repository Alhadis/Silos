// ram holding the test program
module ram(
    input wire [13:0] address,
    input wire [7:0] wdata,
    input wire rw,
    input wire ce,
    output wire [7:0] rdata);

reg [7:0] mem[0:16383];

assign rdata = (ce && rw) ? mem[address] : 8'bz;

always @(posedge rw)
begin
    if (ce)
        mem[address] <= wdata;
end

initial begin
//    $readmemh("cpu6502/tests/functional/test.hexdump", mem);
mem[0] = 8'h00;
mem[1] = 8'h00;
mem[2] = 8'h00;
mem[3] = 8'h00;
mem[4] = 8'h00;
mem[5] = 8'h00;
mem[6] = 8'h00;
mem[7] = 8'h00;
mem[8] = 8'h00;
mem[9] = 8'h00;
mem[10] = 8'h00;
mem[11] = 8'h00;
mem[12] = 8'h00;
mem[13] = 8'h00;
mem[14] = 8'h00;
mem[15] = 8'h00;
mem[16] = 8'h00;
mem[17] = 8'h00;
mem[18] = 8'h00;
mem[19] = 8'h00;
mem[20] = 8'h00;
mem[21] = 8'h00;
mem[22] = 8'h00;
mem[23] = 8'h00;
mem[24] = 8'h00;
mem[25] = 8'h00;
mem[26] = 8'h00;
mem[27] = 8'h00;
mem[28] = 8'h00;
mem[29] = 8'h00;
mem[30] = 8'h00;
mem[31] = 8'h00;
mem[32] = 8'h00;
mem[33] = 8'h00;
mem[34] = 8'h00;
mem[35] = 8'h00;
mem[36] = 8'h00;
mem[37] = 8'h00;
mem[38] = 8'h00;
mem[39] = 8'h00;
mem[40] = 8'h00;
mem[41] = 8'h00;
mem[42] = 8'h00;
mem[43] = 8'h00;
mem[44] = 8'h00;
mem[45] = 8'h00;
mem[46] = 8'h00;
mem[47] = 8'h00;
mem[48] = 8'h00;
mem[49] = 8'h00;
mem[50] = 8'h00;
mem[51] = 8'h00;
mem[52] = 8'h00;
mem[53] = 8'h00;
mem[54] = 8'h00;
mem[55] = 8'h00;
mem[56] = 8'h00;
mem[57] = 8'h00;
mem[58] = 8'h00;
mem[59] = 8'h00;
mem[60] = 8'h00;
mem[61] = 8'h00;
mem[62] = 8'h00;
mem[63] = 8'h00;
mem[64] = 8'h00;
mem[65] = 8'h00;
mem[66] = 8'h00;
mem[67] = 8'h00;
mem[68] = 8'h00;
mem[69] = 8'h00;
mem[70] = 8'h00;
mem[71] = 8'h00;
mem[72] = 8'h00;
mem[73] = 8'h00;
mem[74] = 8'h00;
mem[75] = 8'h00;
mem[76] = 8'h00;
mem[77] = 8'h00;
mem[78] = 8'h00;
mem[79] = 8'h00;
mem[80] = 8'h00;
mem[81] = 8'h00;
mem[82] = 8'h00;
mem[83] = 8'h00;
mem[84] = 8'h00;
mem[85] = 8'h00;
mem[86] = 8'h00;
mem[87] = 8'h00;
mem[88] = 8'h00;
mem[89] = 8'h00;
mem[90] = 8'h00;
mem[91] = 8'h00;
mem[92] = 8'h00;
mem[93] = 8'h00;
mem[94] = 8'h00;
mem[95] = 8'h00;
mem[96] = 8'h00;
mem[97] = 8'h00;
mem[98] = 8'h00;
mem[99] = 8'h00;
mem[100] = 8'h00;
mem[101] = 8'h00;
mem[102] = 8'h00;
mem[103] = 8'h00;
mem[104] = 8'h00;
mem[105] = 8'h00;
mem[106] = 8'h00;
mem[107] = 8'h00;
mem[108] = 8'h00;
mem[109] = 8'h00;
mem[110] = 8'h00;
mem[111] = 8'h00;
mem[112] = 8'h00;
mem[113] = 8'h00;
mem[114] = 8'h00;
mem[115] = 8'h00;
mem[116] = 8'h00;
mem[117] = 8'h00;
mem[118] = 8'h00;
mem[119] = 8'h00;
mem[120] = 8'h00;
mem[121] = 8'h00;
mem[122] = 8'h00;
mem[123] = 8'h00;
mem[124] = 8'h00;
mem[125] = 8'h00;
mem[126] = 8'h00;
mem[127] = 8'h00;
mem[128] = 8'h00;
mem[129] = 8'h00;
mem[130] = 8'h00;
mem[131] = 8'h00;
mem[132] = 8'h00;
mem[133] = 8'h00;
mem[134] = 8'h00;
mem[135] = 8'h00;
mem[136] = 8'h00;
mem[137] = 8'h00;
mem[138] = 8'h00;
mem[139] = 8'h00;
mem[140] = 8'h00;
mem[141] = 8'h00;
mem[142] = 8'h00;
mem[143] = 8'h00;
mem[144] = 8'h00;
mem[145] = 8'h00;
mem[146] = 8'h00;
mem[147] = 8'h00;
mem[148] = 8'h00;
mem[149] = 8'h00;
mem[150] = 8'h00;
mem[151] = 8'h00;
mem[152] = 8'h00;
mem[153] = 8'h00;
mem[154] = 8'h00;
mem[155] = 8'h00;
mem[156] = 8'h00;
mem[157] = 8'h00;
mem[158] = 8'h00;
mem[159] = 8'h00;
mem[160] = 8'h00;
mem[161] = 8'h00;
mem[162] = 8'h00;
mem[163] = 8'h00;
mem[164] = 8'h00;
mem[165] = 8'h00;
mem[166] = 8'h00;
mem[167] = 8'h00;
mem[168] = 8'h00;
mem[169] = 8'h00;
mem[170] = 8'h00;
mem[171] = 8'h00;
mem[172] = 8'h00;
mem[173] = 8'h00;
mem[174] = 8'h00;
mem[175] = 8'h00;
mem[176] = 8'h00;
mem[177] = 8'h00;
mem[178] = 8'h00;
mem[179] = 8'h00;
mem[180] = 8'h00;
mem[181] = 8'h00;
mem[182] = 8'h00;
mem[183] = 8'h00;
mem[184] = 8'h00;
mem[185] = 8'h00;
mem[186] = 8'h00;
mem[187] = 8'h00;
mem[188] = 8'h00;
mem[189] = 8'h00;
mem[190] = 8'h00;
mem[191] = 8'h00;
mem[192] = 8'h00;
mem[193] = 8'h00;
mem[194] = 8'h00;
mem[195] = 8'h00;
mem[196] = 8'h00;
mem[197] = 8'h00;
mem[198] = 8'h00;
mem[199] = 8'h00;
mem[200] = 8'h00;
mem[201] = 8'h00;
mem[202] = 8'h00;
mem[203] = 8'h00;
mem[204] = 8'h00;
mem[205] = 8'h00;
mem[206] = 8'h00;
mem[207] = 8'h00;
mem[208] = 8'h00;
mem[209] = 8'h00;
mem[210] = 8'h00;
mem[211] = 8'h00;
mem[212] = 8'h00;
mem[213] = 8'h00;
mem[214] = 8'h00;
mem[215] = 8'h00;
mem[216] = 8'h00;
mem[217] = 8'h00;
mem[218] = 8'h00;
mem[219] = 8'h00;
mem[220] = 8'h00;
mem[221] = 8'h00;
mem[222] = 8'h00;
mem[223] = 8'h00;
mem[224] = 8'h00;
mem[225] = 8'h00;
mem[226] = 8'h00;
mem[227] = 8'h00;
mem[228] = 8'h00;
mem[229] = 8'h00;
mem[230] = 8'h00;
mem[231] = 8'h00;
mem[232] = 8'h00;
mem[233] = 8'h00;
mem[234] = 8'h00;
mem[235] = 8'h00;
mem[236] = 8'h00;
mem[237] = 8'h00;
mem[238] = 8'h00;
mem[239] = 8'h00;
mem[240] = 8'h00;
mem[241] = 8'h00;
mem[242] = 8'h00;
mem[243] = 8'h00;
mem[244] = 8'h00;
mem[245] = 8'h00;
mem[246] = 8'h00;
mem[247] = 8'h00;
mem[248] = 8'h00;
mem[249] = 8'h00;
mem[250] = 8'h00;
mem[251] = 8'h00;
mem[252] = 8'h00;
mem[253] = 8'h00;
mem[254] = 8'h00;
mem[255] = 8'h00;
mem[256] = 8'h00;
mem[257] = 8'h00;
mem[258] = 8'h00;
mem[259] = 8'h00;
mem[260] = 8'h00;
mem[261] = 8'h00;
mem[262] = 8'h00;
mem[263] = 8'h00;
mem[264] = 8'h00;
mem[265] = 8'h00;
mem[266] = 8'h00;
mem[267] = 8'h00;
mem[268] = 8'h00;
mem[269] = 8'h00;
mem[270] = 8'h00;
mem[271] = 8'h00;
mem[272] = 8'h00;
mem[273] = 8'h00;
mem[274] = 8'h00;
mem[275] = 8'h00;
mem[276] = 8'h00;
mem[277] = 8'h00;
mem[278] = 8'h00;
mem[279] = 8'h00;
mem[280] = 8'h00;
mem[281] = 8'h00;
mem[282] = 8'h00;
mem[283] = 8'h00;
mem[284] = 8'h00;
mem[285] = 8'h00;
mem[286] = 8'h00;
mem[287] = 8'h00;
mem[288] = 8'h00;
mem[289] = 8'h00;
mem[290] = 8'h00;
mem[291] = 8'h00;
mem[292] = 8'h00;
mem[293] = 8'h00;
mem[294] = 8'h00;
mem[295] = 8'h00;
mem[296] = 8'h00;
mem[297] = 8'h00;
mem[298] = 8'h00;
mem[299] = 8'h00;
mem[300] = 8'h00;
mem[301] = 8'h00;
mem[302] = 8'h00;
mem[303] = 8'h00;
mem[304] = 8'h00;
mem[305] = 8'h00;
mem[306] = 8'h00;
mem[307] = 8'h00;
mem[308] = 8'h00;
mem[309] = 8'h00;
mem[310] = 8'h00;
mem[311] = 8'h00;
mem[312] = 8'h00;
mem[313] = 8'h00;
mem[314] = 8'h00;
mem[315] = 8'h00;
mem[316] = 8'h00;
mem[317] = 8'h00;
mem[318] = 8'h00;
mem[319] = 8'h00;
mem[320] = 8'h00;
mem[321] = 8'h00;
mem[322] = 8'h00;
mem[323] = 8'h00;
mem[324] = 8'h00;
mem[325] = 8'h00;
mem[326] = 8'h00;
mem[327] = 8'h00;
mem[328] = 8'h00;
mem[329] = 8'h00;
mem[330] = 8'h00;
mem[331] = 8'h00;
mem[332] = 8'h00;
mem[333] = 8'h00;
mem[334] = 8'h00;
mem[335] = 8'h00;
mem[336] = 8'h00;
mem[337] = 8'h00;
mem[338] = 8'h00;
mem[339] = 8'h00;
mem[340] = 8'h00;
mem[341] = 8'h00;
mem[342] = 8'h00;
mem[343] = 8'h00;
mem[344] = 8'h00;
mem[345] = 8'h00;
mem[346] = 8'h00;
mem[347] = 8'h00;
mem[348] = 8'h00;
mem[349] = 8'h00;
mem[350] = 8'h00;
mem[351] = 8'h00;
mem[352] = 8'h00;
mem[353] = 8'h00;
mem[354] = 8'h00;
mem[355] = 8'h00;
mem[356] = 8'h00;
mem[357] = 8'h00;
mem[358] = 8'h00;
mem[359] = 8'h00;
mem[360] = 8'h00;
mem[361] = 8'h00;
mem[362] = 8'h00;
mem[363] = 8'h00;
mem[364] = 8'h00;
mem[365] = 8'h00;
mem[366] = 8'h00;
mem[367] = 8'h00;
mem[368] = 8'h00;
mem[369] = 8'h00;
mem[370] = 8'h00;
mem[371] = 8'h00;
mem[372] = 8'h00;
mem[373] = 8'h00;
mem[374] = 8'h00;
mem[375] = 8'h00;
mem[376] = 8'h00;
mem[377] = 8'h00;
mem[378] = 8'h00;
mem[379] = 8'h00;
mem[380] = 8'h00;
mem[381] = 8'h00;
mem[382] = 8'h00;
mem[383] = 8'h00;
mem[384] = 8'h00;
mem[385] = 8'h00;
mem[386] = 8'h00;
mem[387] = 8'h00;
mem[388] = 8'h00;
mem[389] = 8'h00;
mem[390] = 8'h00;
mem[391] = 8'h00;
mem[392] = 8'h00;
mem[393] = 8'h00;
mem[394] = 8'h00;
mem[395] = 8'h00;
mem[396] = 8'h00;
mem[397] = 8'h00;
mem[398] = 8'h00;
mem[399] = 8'h00;
mem[400] = 8'h00;
mem[401] = 8'h00;
mem[402] = 8'h00;
mem[403] = 8'h00;
mem[404] = 8'h00;
mem[405] = 8'h00;
mem[406] = 8'h00;
mem[407] = 8'h00;
mem[408] = 8'h00;
mem[409] = 8'h00;
mem[410] = 8'h00;
mem[411] = 8'h00;
mem[412] = 8'h00;
mem[413] = 8'h00;
mem[414] = 8'h00;
mem[415] = 8'h00;
mem[416] = 8'h00;
mem[417] = 8'h00;
mem[418] = 8'h00;
mem[419] = 8'h00;
mem[420] = 8'h00;
mem[421] = 8'h00;
mem[422] = 8'h00;
mem[423] = 8'h00;
mem[424] = 8'h00;
mem[425] = 8'h00;
mem[426] = 8'h00;
mem[427] = 8'h00;
mem[428] = 8'h00;
mem[429] = 8'h00;
mem[430] = 8'h00;
mem[431] = 8'h00;
mem[432] = 8'h00;
mem[433] = 8'h00;
mem[434] = 8'h00;
mem[435] = 8'h00;
mem[436] = 8'h00;
mem[437] = 8'h00;
mem[438] = 8'h00;
mem[439] = 8'h00;
mem[440] = 8'h00;
mem[441] = 8'h00;
mem[442] = 8'h00;
mem[443] = 8'h00;
mem[444] = 8'h00;
mem[445] = 8'h00;
mem[446] = 8'h00;
mem[447] = 8'h00;
mem[448] = 8'h00;
mem[449] = 8'h00;
mem[450] = 8'h00;
mem[451] = 8'h00;
mem[452] = 8'h00;
mem[453] = 8'h00;
mem[454] = 8'h00;
mem[455] = 8'h00;
mem[456] = 8'h00;
mem[457] = 8'h00;
mem[458] = 8'h00;
mem[459] = 8'h00;
mem[460] = 8'h00;
mem[461] = 8'h00;
mem[462] = 8'h00;
mem[463] = 8'h00;
mem[464] = 8'h00;
mem[465] = 8'h00;
mem[466] = 8'h00;
mem[467] = 8'h00;
mem[468] = 8'h00;
mem[469] = 8'h00;
mem[470] = 8'h00;
mem[471] = 8'h00;
mem[472] = 8'h00;
mem[473] = 8'h00;
mem[474] = 8'h00;
mem[475] = 8'h00;
mem[476] = 8'h00;
mem[477] = 8'h00;
mem[478] = 8'h00;
mem[479] = 8'h00;
mem[480] = 8'h00;
mem[481] = 8'h00;
mem[482] = 8'h00;
mem[483] = 8'h00;
mem[484] = 8'h00;
mem[485] = 8'h00;
mem[486] = 8'h00;
mem[487] = 8'h00;
mem[488] = 8'h00;
mem[489] = 8'h00;
mem[490] = 8'h00;
mem[491] = 8'h00;
mem[492] = 8'h00;
mem[493] = 8'h00;
mem[494] = 8'h00;
mem[495] = 8'h00;
mem[496] = 8'h00;
mem[497] = 8'h00;
mem[498] = 8'h00;
mem[499] = 8'h00;
mem[500] = 8'h00;
mem[501] = 8'h00;
mem[502] = 8'h00;
mem[503] = 8'h00;
mem[504] = 8'h00;
mem[505] = 8'h00;
mem[506] = 8'h00;
mem[507] = 8'h00;
mem[508] = 8'h00;
mem[509] = 8'h00;
mem[510] = 8'h00;
mem[511] = 8'h00;
mem[512] = 8'h00;
mem[513] = 8'h00;
mem[514] = 8'h00;
mem[515] = 8'h00;
mem[516] = 8'h00;
mem[517] = 8'h00;
mem[518] = 8'h00;
mem[519] = 8'h00;
mem[520] = 8'h00;
mem[521] = 8'h00;
mem[522] = 8'h00;
mem[523] = 8'h00;
mem[524] = 8'h00;
mem[525] = 8'h00;
mem[526] = 8'h00;
mem[527] = 8'h00;
mem[528] = 8'h00;
mem[529] = 8'h00;
mem[530] = 8'h00;
mem[531] = 8'h00;
mem[532] = 8'h00;
mem[533] = 8'h00;
mem[534] = 8'h00;
mem[535] = 8'h00;
mem[536] = 8'h00;
mem[537] = 8'h00;
mem[538] = 8'h00;
mem[539] = 8'h00;
mem[540] = 8'h00;
mem[541] = 8'h00;
mem[542] = 8'h00;
mem[543] = 8'h00;
mem[544] = 8'h00;
mem[545] = 8'h00;
mem[546] = 8'h00;
mem[547] = 8'h00;
mem[548] = 8'h00;
mem[549] = 8'h00;
mem[550] = 8'h00;
mem[551] = 8'h00;
mem[552] = 8'h00;
mem[553] = 8'h00;
mem[554] = 8'h00;
mem[555] = 8'h00;
mem[556] = 8'h00;
mem[557] = 8'h00;
mem[558] = 8'h00;
mem[559] = 8'h00;
mem[560] = 8'h00;
mem[561] = 8'h00;
mem[562] = 8'h00;
mem[563] = 8'h00;
mem[564] = 8'h00;
mem[565] = 8'h00;
mem[566] = 8'h00;
mem[567] = 8'h00;
mem[568] = 8'h00;
mem[569] = 8'h00;
mem[570] = 8'h00;
mem[571] = 8'h00;
mem[572] = 8'h00;
mem[573] = 8'h00;
mem[574] = 8'h00;
mem[575] = 8'h00;
mem[576] = 8'h00;
mem[577] = 8'h00;
mem[578] = 8'h00;
mem[579] = 8'h00;
mem[580] = 8'h00;
mem[581] = 8'h00;
mem[582] = 8'h00;
mem[583] = 8'h00;
mem[584] = 8'h00;
mem[585] = 8'h00;
mem[586] = 8'h00;
mem[587] = 8'h00;
mem[588] = 8'h00;
mem[589] = 8'h00;
mem[590] = 8'h00;
mem[591] = 8'h00;
mem[592] = 8'h00;
mem[593] = 8'h00;
mem[594] = 8'h00;
mem[595] = 8'h00;
mem[596] = 8'h00;
mem[597] = 8'h00;
mem[598] = 8'h00;
mem[599] = 8'h00;
mem[600] = 8'h00;
mem[601] = 8'h00;
mem[602] = 8'h00;
mem[603] = 8'h00;
mem[604] = 8'h00;
mem[605] = 8'h00;
mem[606] = 8'h00;
mem[607] = 8'h00;
mem[608] = 8'h00;
mem[609] = 8'h00;
mem[610] = 8'h00;
mem[611] = 8'h00;
mem[612] = 8'h00;
mem[613] = 8'h00;
mem[614] = 8'h00;
mem[615] = 8'h00;
mem[616] = 8'h00;
mem[617] = 8'h00;
mem[618] = 8'h00;
mem[619] = 8'h00;
mem[620] = 8'h00;
mem[621] = 8'h00;
mem[622] = 8'h00;
mem[623] = 8'h00;
mem[624] = 8'h00;
mem[625] = 8'h00;
mem[626] = 8'h00;
mem[627] = 8'h00;
mem[628] = 8'h00;
mem[629] = 8'h00;
mem[630] = 8'h00;
mem[631] = 8'h00;
mem[632] = 8'h00;
mem[633] = 8'h00;
mem[634] = 8'h00;
mem[635] = 8'h00;
mem[636] = 8'h00;
mem[637] = 8'h00;
mem[638] = 8'h00;
mem[639] = 8'h00;
mem[640] = 8'h00;
mem[641] = 8'h00;
mem[642] = 8'h00;
mem[643] = 8'h00;
mem[644] = 8'h00;
mem[645] = 8'h00;
mem[646] = 8'h00;
mem[647] = 8'h00;
mem[648] = 8'h00;
mem[649] = 8'h00;
mem[650] = 8'h00;
mem[651] = 8'h00;
mem[652] = 8'h00;
mem[653] = 8'h00;
mem[654] = 8'h00;
mem[655] = 8'h00;
mem[656] = 8'h00;
mem[657] = 8'h00;
mem[658] = 8'h00;
mem[659] = 8'h00;
mem[660] = 8'h00;
mem[661] = 8'h00;
mem[662] = 8'h00;
mem[663] = 8'h00;
mem[664] = 8'h00;
mem[665] = 8'h00;
mem[666] = 8'h00;
mem[667] = 8'h00;
mem[668] = 8'h00;
mem[669] = 8'h00;
mem[670] = 8'h00;
mem[671] = 8'h00;
mem[672] = 8'h00;
mem[673] = 8'h00;
mem[674] = 8'h00;
mem[675] = 8'h00;
mem[676] = 8'h00;
mem[677] = 8'h00;
mem[678] = 8'h00;
mem[679] = 8'h00;
mem[680] = 8'h00;
mem[681] = 8'h00;
mem[682] = 8'h00;
mem[683] = 8'h00;
mem[684] = 8'h00;
mem[685] = 8'h00;
mem[686] = 8'h00;
mem[687] = 8'h00;
mem[688] = 8'h00;
mem[689] = 8'h00;
mem[690] = 8'h00;
mem[691] = 8'h00;
mem[692] = 8'h00;
mem[693] = 8'h00;
mem[694] = 8'h00;
mem[695] = 8'h00;
mem[696] = 8'h00;
mem[697] = 8'h00;
mem[698] = 8'h00;
mem[699] = 8'h00;
mem[700] = 8'h00;
mem[701] = 8'h00;
mem[702] = 8'h00;
mem[703] = 8'h00;
mem[704] = 8'h00;
mem[705] = 8'h00;
mem[706] = 8'h00;
mem[707] = 8'h00;
mem[708] = 8'h00;
mem[709] = 8'h00;
mem[710] = 8'h00;
mem[711] = 8'h00;
mem[712] = 8'h00;
mem[713] = 8'h00;
mem[714] = 8'h00;
mem[715] = 8'h00;
mem[716] = 8'h00;
mem[717] = 8'h00;
mem[718] = 8'h00;
mem[719] = 8'h00;
mem[720] = 8'h00;
mem[721] = 8'h00;
mem[722] = 8'h00;
mem[723] = 8'h00;
mem[724] = 8'h00;
mem[725] = 8'h00;
mem[726] = 8'h00;
mem[727] = 8'h00;
mem[728] = 8'h00;
mem[729] = 8'h00;
mem[730] = 8'h00;
mem[731] = 8'h00;
mem[732] = 8'h00;
mem[733] = 8'h00;
mem[734] = 8'h00;
mem[735] = 8'h00;
mem[736] = 8'h00;
mem[737] = 8'h00;
mem[738] = 8'h00;
mem[739] = 8'h00;
mem[740] = 8'h00;
mem[741] = 8'h00;
mem[742] = 8'h00;
mem[743] = 8'h00;
mem[744] = 8'h00;
mem[745] = 8'h00;
mem[746] = 8'h00;
mem[747] = 8'h00;
mem[748] = 8'h00;
mem[749] = 8'h00;
mem[750] = 8'h00;
mem[751] = 8'h00;
mem[752] = 8'h00;
mem[753] = 8'h00;
mem[754] = 8'h00;
mem[755] = 8'h00;
mem[756] = 8'h00;
mem[757] = 8'h00;
mem[758] = 8'h00;
mem[759] = 8'h00;
mem[760] = 8'h00;
mem[761] = 8'h00;
mem[762] = 8'h00;
mem[763] = 8'h00;
mem[764] = 8'h00;
mem[765] = 8'h00;
mem[766] = 8'h00;
mem[767] = 8'h00;
mem[768] = 8'h00;
mem[769] = 8'h00;
mem[770] = 8'h00;
mem[771] = 8'h00;
mem[772] = 8'h00;
mem[773] = 8'h00;
mem[774] = 8'h00;
mem[775] = 8'h00;
mem[776] = 8'h00;
mem[777] = 8'h00;
mem[778] = 8'h00;
mem[779] = 8'h00;
mem[780] = 8'h00;
mem[781] = 8'h00;
mem[782] = 8'h00;
mem[783] = 8'h00;
mem[784] = 8'h00;
mem[785] = 8'h00;
mem[786] = 8'h00;
mem[787] = 8'h00;
mem[788] = 8'h00;
mem[789] = 8'h00;
mem[790] = 8'h00;
mem[791] = 8'h00;
mem[792] = 8'h00;
mem[793] = 8'h00;
mem[794] = 8'h00;
mem[795] = 8'h00;
mem[796] = 8'h00;
mem[797] = 8'h00;
mem[798] = 8'h00;
mem[799] = 8'h00;
mem[800] = 8'h00;
mem[801] = 8'h00;
mem[802] = 8'h00;
mem[803] = 8'h00;
mem[804] = 8'h00;
mem[805] = 8'h00;
mem[806] = 8'h00;
mem[807] = 8'h00;
mem[808] = 8'h00;
mem[809] = 8'h00;
mem[810] = 8'h00;
mem[811] = 8'h00;
mem[812] = 8'h00;
mem[813] = 8'h00;
mem[814] = 8'h00;
mem[815] = 8'h00;
mem[816] = 8'h00;
mem[817] = 8'h00;
mem[818] = 8'h00;
mem[819] = 8'h00;
mem[820] = 8'h00;
mem[821] = 8'h00;
mem[822] = 8'h00;
mem[823] = 8'h00;
mem[824] = 8'h00;
mem[825] = 8'h00;
mem[826] = 8'h00;
mem[827] = 8'h00;
mem[828] = 8'h00;
mem[829] = 8'h00;
mem[830] = 8'h00;
mem[831] = 8'h00;
mem[832] = 8'h00;
mem[833] = 8'h00;
mem[834] = 8'h00;
mem[835] = 8'h00;
mem[836] = 8'h00;
mem[837] = 8'h00;
mem[838] = 8'h00;
mem[839] = 8'h00;
mem[840] = 8'h00;
mem[841] = 8'h00;
mem[842] = 8'h00;
mem[843] = 8'h00;
mem[844] = 8'h00;
mem[845] = 8'h00;
mem[846] = 8'h00;
mem[847] = 8'h00;
mem[848] = 8'h00;
mem[849] = 8'h00;
mem[850] = 8'h00;
mem[851] = 8'h00;
mem[852] = 8'h00;
mem[853] = 8'h00;
mem[854] = 8'h00;
mem[855] = 8'h00;
mem[856] = 8'h00;
mem[857] = 8'h00;
mem[858] = 8'h00;
mem[859] = 8'h00;
mem[860] = 8'h00;
mem[861] = 8'h00;
mem[862] = 8'h00;
mem[863] = 8'h00;
mem[864] = 8'h00;
mem[865] = 8'h00;
mem[866] = 8'h00;
mem[867] = 8'h00;
mem[868] = 8'h00;
mem[869] = 8'h00;
mem[870] = 8'h00;
mem[871] = 8'h00;
mem[872] = 8'h00;
mem[873] = 8'h00;
mem[874] = 8'h00;
mem[875] = 8'h00;
mem[876] = 8'h00;
mem[877] = 8'h00;
mem[878] = 8'h00;
mem[879] = 8'h00;
mem[880] = 8'h00;
mem[881] = 8'h00;
mem[882] = 8'h00;
mem[883] = 8'h00;
mem[884] = 8'h00;
mem[885] = 8'h00;
mem[886] = 8'h00;
mem[887] = 8'h00;
mem[888] = 8'h00;
mem[889] = 8'h00;
mem[890] = 8'h00;
mem[891] = 8'h00;
mem[892] = 8'h00;
mem[893] = 8'h00;
mem[894] = 8'h00;
mem[895] = 8'h00;
mem[896] = 8'h00;
mem[897] = 8'h00;
mem[898] = 8'h00;
mem[899] = 8'h00;
mem[900] = 8'h00;
mem[901] = 8'h00;
mem[902] = 8'h00;
mem[903] = 8'h00;
mem[904] = 8'h00;
mem[905] = 8'h00;
mem[906] = 8'h00;
mem[907] = 8'h00;
mem[908] = 8'h00;
mem[909] = 8'h00;
mem[910] = 8'h00;
mem[911] = 8'h00;
mem[912] = 8'h00;
mem[913] = 8'h00;
mem[914] = 8'h00;
mem[915] = 8'h00;
mem[916] = 8'h00;
mem[917] = 8'h00;
mem[918] = 8'h00;
mem[919] = 8'h00;
mem[920] = 8'h00;
mem[921] = 8'h00;
mem[922] = 8'h00;
mem[923] = 8'h00;
mem[924] = 8'h00;
mem[925] = 8'h00;
mem[926] = 8'h00;
mem[927] = 8'h00;
mem[928] = 8'h00;
mem[929] = 8'h00;
mem[930] = 8'h00;
mem[931] = 8'h00;
mem[932] = 8'h00;
mem[933] = 8'h00;
mem[934] = 8'h00;
mem[935] = 8'h00;
mem[936] = 8'h00;
mem[937] = 8'h00;
mem[938] = 8'h00;
mem[939] = 8'h00;
mem[940] = 8'h00;
mem[941] = 8'h00;
mem[942] = 8'h00;
mem[943] = 8'h00;
mem[944] = 8'h00;
mem[945] = 8'h00;
mem[946] = 8'h00;
mem[947] = 8'h00;
mem[948] = 8'h00;
mem[949] = 8'h00;
mem[950] = 8'h00;
mem[951] = 8'h00;
mem[952] = 8'h00;
mem[953] = 8'h00;
mem[954] = 8'h00;
mem[955] = 8'h00;
mem[956] = 8'h00;
mem[957] = 8'h00;
mem[958] = 8'h00;
mem[959] = 8'h00;
mem[960] = 8'h00;
mem[961] = 8'h00;
mem[962] = 8'h00;
mem[963] = 8'h00;
mem[964] = 8'h00;
mem[965] = 8'h00;
mem[966] = 8'h00;
mem[967] = 8'h00;
mem[968] = 8'h00;
mem[969] = 8'h00;
mem[970] = 8'h00;
mem[971] = 8'h00;
mem[972] = 8'h00;
mem[973] = 8'h00;
mem[974] = 8'h00;
mem[975] = 8'h00;
mem[976] = 8'h00;
mem[977] = 8'h00;
mem[978] = 8'h00;
mem[979] = 8'h00;
mem[980] = 8'h00;
mem[981] = 8'h00;
mem[982] = 8'h00;
mem[983] = 8'h00;
mem[984] = 8'h00;
mem[985] = 8'h00;
mem[986] = 8'h00;
mem[987] = 8'h00;
mem[988] = 8'h00;
mem[989] = 8'h00;
mem[990] = 8'h00;
mem[991] = 8'h00;
mem[992] = 8'h00;
mem[993] = 8'h00;
mem[994] = 8'h00;
mem[995] = 8'h00;
mem[996] = 8'h00;
mem[997] = 8'h00;
mem[998] = 8'h00;
mem[999] = 8'h00;
mem[1000] = 8'h00;
mem[1001] = 8'h00;
mem[1002] = 8'h00;
mem[1003] = 8'h00;
mem[1004] = 8'h00;
mem[1005] = 8'h00;
mem[1006] = 8'h00;
mem[1007] = 8'h00;
mem[1008] = 8'h00;
mem[1009] = 8'h00;
mem[1010] = 8'h00;
mem[1011] = 8'h00;
mem[1012] = 8'h00;
mem[1013] = 8'h00;
mem[1014] = 8'h00;
mem[1015] = 8'h00;
mem[1016] = 8'h00;
mem[1017] = 8'h00;
mem[1018] = 8'h00;
mem[1019] = 8'h00;
mem[1020] = 8'h00;
mem[1021] = 8'h00;
mem[1022] = 8'h00;
mem[1023] = 8'h00;
mem[1024] = 8'hd8;
mem[1025] = 8'ha2;
mem[1026] = 8'hff;
mem[1027] = 8'h9a;
mem[1028] = 8'ha9;
mem[1029] = 8'h00;
mem[1030] = 8'h8d;
mem[1031] = 8'h00;
mem[1032] = 8'h02;
mem[1033] = 8'ha2;
mem[1034] = 8'h05;
mem[1035] = 8'h4c;
mem[1036] = 8'h33;
mem[1037] = 8'h04;
mem[1038] = 8'ha0;
mem[1039] = 8'h05;
mem[1040] = 8'hd0;
mem[1041] = 8'h08;
mem[1042] = 8'h4c;
mem[1043] = 8'h12;
mem[1044] = 8'h04;
mem[1045] = 8'h88;
mem[1046] = 8'h88;
mem[1047] = 8'h88;
mem[1048] = 8'h88;
mem[1049] = 8'h88;
mem[1050] = 8'h88;
mem[1051] = 8'h88;
mem[1052] = 8'h88;
mem[1053] = 8'h88;
mem[1054] = 8'h88;
mem[1055] = 8'hf0;
mem[1056] = 8'h17;
mem[1057] = 8'h4c;
mem[1058] = 8'h21;
mem[1059] = 8'h04;
mem[1060] = 8'hca;
mem[1061] = 8'hca;
mem[1062] = 8'hca;
mem[1063] = 8'hca;
mem[1064] = 8'hca;
mem[1065] = 8'hca;
mem[1066] = 8'hca;
mem[1067] = 8'hca;
mem[1068] = 8'hca;
mem[1069] = 8'hca;
mem[1070] = 8'hf0;
mem[1071] = 8'hde;
mem[1072] = 8'h4c;
mem[1073] = 8'h30;
mem[1074] = 8'h04;
mem[1075] = 8'hd0;
mem[1076] = 8'hf4;
mem[1077] = 8'h4c;
mem[1078] = 8'h35;
mem[1079] = 8'h04;
mem[1080] = 8'ha2;
mem[1081] = 8'h46;
mem[1082] = 8'hbd;
mem[1083] = 8'hd8;
mem[1084] = 8'h38;
mem[1085] = 8'h95;
mem[1086] = 8'h13;
mem[1087] = 8'hca;
mem[1088] = 8'h10;
mem[1089] = 8'hf8;
mem[1090] = 8'ha2;
mem[1091] = 8'h61;
mem[1092] = 8'hbd;
mem[1093] = 8'h1f;
mem[1094] = 8'h39;
mem[1095] = 8'h9d;
mem[1096] = 8'h08;
mem[1097] = 8'h02;
mem[1098] = 8'hca;
mem[1099] = 8'h10;
mem[1100] = 8'hf7;
mem[1101] = 8'ha2;
mem[1102] = 8'h05;
mem[1103] = 8'hbd;
mem[1104] = 8'h81;
mem[1105] = 8'h39;
mem[1106] = 8'h9d;
mem[1107] = 8'hfa;
mem[1108] = 8'hff;
mem[1109] = 8'hca;
mem[1110] = 8'h10;
mem[1111] = 8'hf7;
mem[1112] = 8'had;
mem[1113] = 8'h00;
mem[1114] = 8'h02;
mem[1115] = 8'hc9;
mem[1116] = 8'h00;
mem[1117] = 8'hd0;
mem[1118] = 8'hfe;
mem[1119] = 8'ha9;
mem[1120] = 8'h01;
mem[1121] = 8'h8d;
mem[1122] = 8'h00;
mem[1123] = 8'h02;
mem[1124] = 8'ha0;
mem[1125] = 8'hfe;
mem[1126] = 8'h88;
mem[1127] = 8'h98;
mem[1128] = 8'haa;
mem[1129] = 8'h10;
mem[1130] = 8'h08;
mem[1131] = 8'h18;
mem[1132] = 8'h69;
mem[1133] = 8'h02;
mem[1134] = 8'hea;
mem[1135] = 8'hea;
mem[1136] = 8'hea;
mem[1137] = 8'hea;
mem[1138] = 8'hea;
mem[1139] = 8'hea;
mem[1140] = 8'hea;
mem[1141] = 8'hea;
mem[1142] = 8'hea;
mem[1143] = 8'hea;
mem[1144] = 8'h49;
mem[1145] = 8'h7f;
mem[1146] = 8'h8d;
mem[1147] = 8'h06;
mem[1148] = 8'h05;
mem[1149] = 8'ha9;
mem[1150] = 8'h00;
mem[1151] = 8'h4c;
mem[1152] = 8'h05;
mem[1153] = 8'h05;
mem[1154] = 8'hca;
mem[1155] = 8'hca;
mem[1156] = 8'hca;
mem[1157] = 8'hca;
mem[1158] = 8'hca;
mem[1159] = 8'hca;
mem[1160] = 8'hca;
mem[1161] = 8'hca;
mem[1162] = 8'hca;
mem[1163] = 8'hca;
mem[1164] = 8'hca;
mem[1165] = 8'hca;
mem[1166] = 8'hca;
mem[1167] = 8'hca;
mem[1168] = 8'hca;
mem[1169] = 8'hca;
mem[1170] = 8'hca;
mem[1171] = 8'hca;
mem[1172] = 8'hca;
mem[1173] = 8'hca;
mem[1174] = 8'hca;
mem[1175] = 8'hca;
mem[1176] = 8'hca;
mem[1177] = 8'hca;
mem[1178] = 8'hca;
mem[1179] = 8'hca;
mem[1180] = 8'hca;
mem[1181] = 8'hca;
mem[1182] = 8'hca;
mem[1183] = 8'hca;
mem[1184] = 8'hca;
mem[1185] = 8'hca;
mem[1186] = 8'hca;
mem[1187] = 8'hca;
mem[1188] = 8'hca;
mem[1189] = 8'hca;
mem[1190] = 8'hca;
mem[1191] = 8'hca;
mem[1192] = 8'hca;
mem[1193] = 8'hca;
mem[1194] = 8'hca;
mem[1195] = 8'hca;
mem[1196] = 8'hca;
mem[1197] = 8'hca;
mem[1198] = 8'hca;
mem[1199] = 8'hca;
mem[1200] = 8'hca;
mem[1201] = 8'hca;
mem[1202] = 8'hca;
mem[1203] = 8'hca;
mem[1204] = 8'hca;
mem[1205] = 8'hca;
mem[1206] = 8'hca;
mem[1207] = 8'hca;
mem[1208] = 8'hca;
mem[1209] = 8'hca;
mem[1210] = 8'hca;
mem[1211] = 8'hca;
mem[1212] = 8'hca;
mem[1213] = 8'hca;
mem[1214] = 8'hca;
mem[1215] = 8'hca;
mem[1216] = 8'hca;
mem[1217] = 8'hca;
mem[1218] = 8'hca;
mem[1219] = 8'hca;
mem[1220] = 8'hca;
mem[1221] = 8'hca;
mem[1222] = 8'hca;
mem[1223] = 8'hca;
mem[1224] = 8'hca;
mem[1225] = 8'hca;
mem[1226] = 8'hca;
mem[1227] = 8'hca;
mem[1228] = 8'hca;
mem[1229] = 8'hca;
mem[1230] = 8'hca;
mem[1231] = 8'hca;
mem[1232] = 8'hca;
mem[1233] = 8'hca;
mem[1234] = 8'hca;
mem[1235] = 8'hca;
mem[1236] = 8'hca;
mem[1237] = 8'hca;
mem[1238] = 8'hca;
mem[1239] = 8'hca;
mem[1240] = 8'hca;
mem[1241] = 8'hca;
mem[1242] = 8'hca;
mem[1243] = 8'hca;
mem[1244] = 8'hca;
mem[1245] = 8'hca;
mem[1246] = 8'hca;
mem[1247] = 8'hca;
mem[1248] = 8'hca;
mem[1249] = 8'hca;
mem[1250] = 8'hca;
mem[1251] = 8'hca;
mem[1252] = 8'hca;
mem[1253] = 8'hca;
mem[1254] = 8'hca;
mem[1255] = 8'hca;
mem[1256] = 8'hca;
mem[1257] = 8'hca;
mem[1258] = 8'hca;
mem[1259] = 8'hca;
mem[1260] = 8'hca;
mem[1261] = 8'hca;
mem[1262] = 8'hca;
mem[1263] = 8'hca;
mem[1264] = 8'hca;
mem[1265] = 8'hca;
mem[1266] = 8'hca;
mem[1267] = 8'hca;
mem[1268] = 8'hca;
mem[1269] = 8'hca;
mem[1270] = 8'hca;
mem[1271] = 8'hca;
mem[1272] = 8'hca;
mem[1273] = 8'hca;
mem[1274] = 8'hca;
mem[1275] = 8'hca;
mem[1276] = 8'hca;
mem[1277] = 8'hca;
mem[1278] = 8'hca;
mem[1279] = 8'hca;
mem[1280] = 8'hca;
mem[1281] = 8'hca;
mem[1282] = 8'hca;
mem[1283] = 8'hca;
mem[1284] = 8'hca;
mem[1285] = 8'hf0;
mem[1286] = 8'h3e;
mem[1287] = 8'hca;
mem[1288] = 8'hca;
mem[1289] = 8'hca;
mem[1290] = 8'hca;
mem[1291] = 8'hca;
mem[1292] = 8'hca;
mem[1293] = 8'hca;
mem[1294] = 8'hca;
mem[1295] = 8'hca;
mem[1296] = 8'hca;
mem[1297] = 8'hca;
mem[1298] = 8'hca;
mem[1299] = 8'hca;
mem[1300] = 8'hca;
mem[1301] = 8'hca;
mem[1302] = 8'hca;
mem[1303] = 8'hca;
mem[1304] = 8'hca;
mem[1305] = 8'hca;
mem[1306] = 8'hca;
mem[1307] = 8'hca;
mem[1308] = 8'hca;
mem[1309] = 8'hca;
mem[1310] = 8'hca;
mem[1311] = 8'hca;
mem[1312] = 8'hca;
mem[1313] = 8'hca;
mem[1314] = 8'hca;
mem[1315] = 8'hca;
mem[1316] = 8'hca;
mem[1317] = 8'hca;
mem[1318] = 8'hca;
mem[1319] = 8'hca;
mem[1320] = 8'hca;
mem[1321] = 8'hca;
mem[1322] = 8'hca;
mem[1323] = 8'hca;
mem[1324] = 8'hca;
mem[1325] = 8'hca;
mem[1326] = 8'hca;
mem[1327] = 8'hca;
mem[1328] = 8'hca;
mem[1329] = 8'hca;
mem[1330] = 8'hca;
mem[1331] = 8'hca;
mem[1332] = 8'hca;
mem[1333] = 8'hca;
mem[1334] = 8'hca;
mem[1335] = 8'hca;
mem[1336] = 8'hca;
mem[1337] = 8'hca;
mem[1338] = 8'hca;
mem[1339] = 8'hca;
mem[1340] = 8'hca;
mem[1341] = 8'hca;
mem[1342] = 8'hca;
mem[1343] = 8'hca;
mem[1344] = 8'hca;
mem[1345] = 8'hca;
mem[1346] = 8'hca;
mem[1347] = 8'hca;
mem[1348] = 8'hca;
mem[1349] = 8'hca;
mem[1350] = 8'hca;
mem[1351] = 8'hca;
mem[1352] = 8'hca;
mem[1353] = 8'hca;
mem[1354] = 8'hca;
mem[1355] = 8'hca;
mem[1356] = 8'hca;
mem[1357] = 8'hca;
mem[1358] = 8'hca;
mem[1359] = 8'hca;
mem[1360] = 8'hca;
mem[1361] = 8'hca;
mem[1362] = 8'hca;
mem[1363] = 8'hca;
mem[1364] = 8'hca;
mem[1365] = 8'hca;
mem[1366] = 8'hca;
mem[1367] = 8'hca;
mem[1368] = 8'hca;
mem[1369] = 8'hca;
mem[1370] = 8'hca;
mem[1371] = 8'hca;
mem[1372] = 8'hca;
mem[1373] = 8'hca;
mem[1374] = 8'hca;
mem[1375] = 8'hca;
mem[1376] = 8'hca;
mem[1377] = 8'hca;
mem[1378] = 8'hca;
mem[1379] = 8'hca;
mem[1380] = 8'hca;
mem[1381] = 8'hca;
mem[1382] = 8'hca;
mem[1383] = 8'hca;
mem[1384] = 8'hca;
mem[1385] = 8'hca;
mem[1386] = 8'hca;
mem[1387] = 8'hca;
mem[1388] = 8'hca;
mem[1389] = 8'hca;
mem[1390] = 8'hca;
mem[1391] = 8'hca;
mem[1392] = 8'hca;
mem[1393] = 8'hca;
mem[1394] = 8'hca;
mem[1395] = 8'hca;
mem[1396] = 8'hca;
mem[1397] = 8'hca;
mem[1398] = 8'hca;
mem[1399] = 8'hca;
mem[1400] = 8'hca;
mem[1401] = 8'hca;
mem[1402] = 8'hca;
mem[1403] = 8'hca;
mem[1404] = 8'hca;
mem[1405] = 8'hca;
mem[1406] = 8'hca;
mem[1407] = 8'hca;
mem[1408] = 8'hca;
mem[1409] = 8'hca;
mem[1410] = 8'hca;
mem[1411] = 8'hca;
mem[1412] = 8'hca;
mem[1413] = 8'hca;
mem[1414] = 8'hea;
mem[1415] = 8'hea;
mem[1416] = 8'hea;
mem[1417] = 8'hea;
mem[1418] = 8'hea;
mem[1419] = 8'hf0;
mem[1420] = 8'h08;
mem[1421] = 8'h4c;
mem[1422] = 8'h8d;
mem[1423] = 8'h05;
mem[1424] = 8'hea;
mem[1425] = 8'hea;
mem[1426] = 8'hea;
mem[1427] = 8'hea;
mem[1428] = 8'hea;
mem[1429] = 8'hea;
mem[1430] = 8'hea;
mem[1431] = 8'hea;
mem[1432] = 8'hea;
mem[1433] = 8'hea;
mem[1434] = 8'hc0;
mem[1435] = 8'h00;
mem[1436] = 8'hf0;
mem[1437] = 8'h03;
mem[1438] = 8'h4c;
mem[1439] = 8'h66;
mem[1440] = 8'h04;
mem[1441] = 8'had;
mem[1442] = 8'h00;
mem[1443] = 8'h02;
mem[1444] = 8'hc9;
mem[1445] = 8'h01;
mem[1446] = 8'hd0;
mem[1447] = 8'hfe;
mem[1448] = 8'ha9;
mem[1449] = 8'h02;
mem[1450] = 8'h8d;
mem[1451] = 8'h00;
mem[1452] = 8'h02;
mem[1453] = 8'hc0;
mem[1454] = 8'h01;
mem[1455] = 8'hd0;
mem[1456] = 8'h03;
mem[1457] = 8'h4c;
mem[1458] = 8'hb1;
mem[1459] = 8'h05;
mem[1460] = 8'ha9;
mem[1461] = 8'h00;
mem[1462] = 8'hc9;
mem[1463] = 8'h00;
mem[1464] = 8'hd0;
mem[1465] = 8'hfe;
mem[1466] = 8'h90;
mem[1467] = 8'hfe;
mem[1468] = 8'h30;
mem[1469] = 8'hfe;
mem[1470] = 8'hc9;
mem[1471] = 8'h01;
mem[1472] = 8'hf0;
mem[1473] = 8'hfe;
mem[1474] = 8'hb0;
mem[1475] = 8'hfe;
mem[1476] = 8'h10;
mem[1477] = 8'hfe;
mem[1478] = 8'haa;
mem[1479] = 8'he0;
mem[1480] = 8'h00;
mem[1481] = 8'hd0;
mem[1482] = 8'hfe;
mem[1483] = 8'h90;
mem[1484] = 8'hfe;
mem[1485] = 8'h30;
mem[1486] = 8'hfe;
mem[1487] = 8'he0;
mem[1488] = 8'h01;
mem[1489] = 8'hf0;
mem[1490] = 8'hfe;
mem[1491] = 8'hb0;
mem[1492] = 8'hfe;
mem[1493] = 8'h10;
mem[1494] = 8'hfe;
mem[1495] = 8'ha8;
mem[1496] = 8'hc0;
mem[1497] = 8'h00;
mem[1498] = 8'hd0;
mem[1499] = 8'hfe;
mem[1500] = 8'h90;
mem[1501] = 8'hfe;
mem[1502] = 8'h30;
mem[1503] = 8'hfe;
mem[1504] = 8'hc0;
mem[1505] = 8'h01;
mem[1506] = 8'hf0;
mem[1507] = 8'hfe;
mem[1508] = 8'hb0;
mem[1509] = 8'hfe;
mem[1510] = 8'h10;
mem[1511] = 8'hfe;
mem[1512] = 8'had;
mem[1513] = 8'h00;
mem[1514] = 8'h02;
mem[1515] = 8'hc9;
mem[1516] = 8'h02;
mem[1517] = 8'hd0;
mem[1518] = 8'hfe;
mem[1519] = 8'ha9;
mem[1520] = 8'h03;
mem[1521] = 8'h8d;
mem[1522] = 8'h00;
mem[1523] = 8'h02;
mem[1524] = 8'ha2;
mem[1525] = 8'hff;
mem[1526] = 8'h9a;
mem[1527] = 8'ha9;
mem[1528] = 8'h55;
mem[1529] = 8'h48;
mem[1530] = 8'ha9;
mem[1531] = 8'haa;
mem[1532] = 8'h48;
mem[1533] = 8'hcd;
mem[1534] = 8'hfe;
mem[1535] = 8'h01;
mem[1536] = 8'hd0;
mem[1537] = 8'hfe;
mem[1538] = 8'hba;
mem[1539] = 8'h8a;
mem[1540] = 8'hc9;
mem[1541] = 8'hfd;
mem[1542] = 8'hd0;
mem[1543] = 8'hfe;
mem[1544] = 8'h68;
mem[1545] = 8'hc9;
mem[1546] = 8'haa;
mem[1547] = 8'hd0;
mem[1548] = 8'hfe;
mem[1549] = 8'h68;
mem[1550] = 8'hc9;
mem[1551] = 8'h55;
mem[1552] = 8'hd0;
mem[1553] = 8'hfe;
mem[1554] = 8'hcd;
mem[1555] = 8'hff;
mem[1556] = 8'h01;
mem[1557] = 8'hd0;
mem[1558] = 8'hfe;
mem[1559] = 8'hba;
mem[1560] = 8'he0;
mem[1561] = 8'hff;
mem[1562] = 8'hd0;
mem[1563] = 8'hfe;
mem[1564] = 8'had;
mem[1565] = 8'h00;
mem[1566] = 8'h02;
mem[1567] = 8'hc9;
mem[1568] = 8'h03;
mem[1569] = 8'hd0;
mem[1570] = 8'hfe;
mem[1571] = 8'ha9;
mem[1572] = 8'h04;
mem[1573] = 8'h8d;
mem[1574] = 8'h00;
mem[1575] = 8'h02;
mem[1576] = 8'ha9;
mem[1577] = 8'hff;
mem[1578] = 8'h48;
mem[1579] = 8'h28;
mem[1580] = 8'h10;
mem[1581] = 8'h1a;
mem[1582] = 8'h50;
mem[1583] = 8'h1b;
mem[1584] = 8'h90;
mem[1585] = 8'h1c;
mem[1586] = 8'hd0;
mem[1587] = 8'h1d;
mem[1588] = 8'h30;
mem[1589] = 8'h03;
mem[1590] = 8'h4c;
mem[1591] = 8'h36;
mem[1592] = 8'h06;
mem[1593] = 8'h70;
mem[1594] = 8'h03;
mem[1595] = 8'h4c;
mem[1596] = 8'h3b;
mem[1597] = 8'h06;
mem[1598] = 8'hb0;
mem[1599] = 8'h03;
mem[1600] = 8'h4c;
mem[1601] = 8'h40;
mem[1602] = 8'h06;
mem[1603] = 8'hf0;
mem[1604] = 8'h0f;
mem[1605] = 8'h4c;
mem[1606] = 8'h45;
mem[1607] = 8'h06;
mem[1608] = 8'h4c;
mem[1609] = 8'h48;
mem[1610] = 8'h06;
mem[1611] = 8'h4c;
mem[1612] = 8'h4b;
mem[1613] = 8'h06;
mem[1614] = 8'h4c;
mem[1615] = 8'h4e;
mem[1616] = 8'h06;
mem[1617] = 8'h4c;
mem[1618] = 8'h51;
mem[1619] = 8'h06;
mem[1620] = 8'h08;
mem[1621] = 8'hba;
mem[1622] = 8'he0;
mem[1623] = 8'hfe;
mem[1624] = 8'hd0;
mem[1625] = 8'hfe;
mem[1626] = 8'h68;
mem[1627] = 8'h09;
mem[1628] = 8'h08;
mem[1629] = 8'hc9;
mem[1630] = 8'hff;
mem[1631] = 8'hd0;
mem[1632] = 8'hfe;
mem[1633] = 8'hba;
mem[1634] = 8'he0;
mem[1635] = 8'hff;
mem[1636] = 8'hd0;
mem[1637] = 8'hfe;
mem[1638] = 8'ha9;
mem[1639] = 8'h00;
mem[1640] = 8'h48;
mem[1641] = 8'h28;
mem[1642] = 8'h30;
mem[1643] = 8'h1a;
mem[1644] = 8'h70;
mem[1645] = 8'h1b;
mem[1646] = 8'hb0;
mem[1647] = 8'h1c;
mem[1648] = 8'hf0;
mem[1649] = 8'h1d;
mem[1650] = 8'h10;
mem[1651] = 8'h03;
mem[1652] = 8'h4c;
mem[1653] = 8'h74;
mem[1654] = 8'h06;
mem[1655] = 8'h50;
mem[1656] = 8'h03;
mem[1657] = 8'h4c;
mem[1658] = 8'h79;
mem[1659] = 8'h06;
mem[1660] = 8'h90;
mem[1661] = 8'h03;
mem[1662] = 8'h4c;
mem[1663] = 8'h7e;
mem[1664] = 8'h06;
mem[1665] = 8'hd0;
mem[1666] = 8'h0f;
mem[1667] = 8'h4c;
mem[1668] = 8'h83;
mem[1669] = 8'h06;
mem[1670] = 8'h4c;
mem[1671] = 8'h86;
mem[1672] = 8'h06;
mem[1673] = 8'h4c;
mem[1674] = 8'h89;
mem[1675] = 8'h06;
mem[1676] = 8'h4c;
mem[1677] = 8'h8c;
mem[1678] = 8'h06;
mem[1679] = 8'h4c;
mem[1680] = 8'h8f;
mem[1681] = 8'h06;
mem[1682] = 8'h08;
mem[1683] = 8'h68;
mem[1684] = 8'h09;
mem[1685] = 8'h08;
mem[1686] = 8'hc9;
mem[1687] = 8'h38;
mem[1688] = 8'hd0;
mem[1689] = 8'hfe;
mem[1690] = 8'ha9;
mem[1691] = 8'h02;
mem[1692] = 8'h48;
mem[1693] = 8'h28;
mem[1694] = 8'hd0;
mem[1695] = 8'h02;
mem[1696] = 8'hf0;
mem[1697] = 8'h03;
mem[1698] = 8'h4c;
mem[1699] = 8'ha2;
mem[1700] = 8'h06;
mem[1701] = 8'hb0;
mem[1702] = 8'h02;
mem[1703] = 8'h90;
mem[1704] = 8'h03;
mem[1705] = 8'h4c;
mem[1706] = 8'ha9;
mem[1707] = 8'h06;
mem[1708] = 8'h30;
mem[1709] = 8'h02;
mem[1710] = 8'h10;
mem[1711] = 8'h03;
mem[1712] = 8'h4c;
mem[1713] = 8'hb0;
mem[1714] = 8'h06;
mem[1715] = 8'h70;
mem[1716] = 8'h02;
mem[1717] = 8'h50;
mem[1718] = 8'h03;
mem[1719] = 8'h4c;
mem[1720] = 8'hb7;
mem[1721] = 8'h06;
mem[1722] = 8'ha9;
mem[1723] = 8'h01;
mem[1724] = 8'h48;
mem[1725] = 8'h28;
mem[1726] = 8'hf0;
mem[1727] = 8'h02;
mem[1728] = 8'hd0;
mem[1729] = 8'h03;
mem[1730] = 8'h4c;
mem[1731] = 8'hc2;
mem[1732] = 8'h06;
mem[1733] = 8'h90;
mem[1734] = 8'h02;
mem[1735] = 8'hb0;
mem[1736] = 8'h03;
mem[1737] = 8'h4c;
mem[1738] = 8'hc9;
mem[1739] = 8'h06;
mem[1740] = 8'h30;
mem[1741] = 8'h02;
mem[1742] = 8'h10;
mem[1743] = 8'h03;
mem[1744] = 8'h4c;
mem[1745] = 8'hd0;
mem[1746] = 8'h06;
mem[1747] = 8'h70;
mem[1748] = 8'h02;
mem[1749] = 8'h50;
mem[1750] = 8'h03;
mem[1751] = 8'h4c;
mem[1752] = 8'hd7;
mem[1753] = 8'h06;
mem[1754] = 8'ha9;
mem[1755] = 8'h80;
mem[1756] = 8'h48;
mem[1757] = 8'h28;
mem[1758] = 8'hf0;
mem[1759] = 8'h02;
mem[1760] = 8'hd0;
mem[1761] = 8'h03;
mem[1762] = 8'h4c;
mem[1763] = 8'he2;
mem[1764] = 8'h06;
mem[1765] = 8'hb0;
mem[1766] = 8'h02;
mem[1767] = 8'h90;
mem[1768] = 8'h03;
mem[1769] = 8'h4c;
mem[1770] = 8'he9;
mem[1771] = 8'h06;
mem[1772] = 8'h10;
mem[1773] = 8'h02;
mem[1774] = 8'h30;
mem[1775] = 8'h03;
mem[1776] = 8'h4c;
mem[1777] = 8'hf0;
mem[1778] = 8'h06;
mem[1779] = 8'h70;
mem[1780] = 8'h02;
mem[1781] = 8'h50;
mem[1782] = 8'h03;
mem[1783] = 8'h4c;
mem[1784] = 8'hf7;
mem[1785] = 8'h06;
mem[1786] = 8'ha9;
mem[1787] = 8'h40;
mem[1788] = 8'h48;
mem[1789] = 8'h28;
mem[1790] = 8'hf0;
mem[1791] = 8'h02;
mem[1792] = 8'hd0;
mem[1793] = 8'h03;
mem[1794] = 8'h4c;
mem[1795] = 8'h02;
mem[1796] = 8'h07;
mem[1797] = 8'hb0;
mem[1798] = 8'h02;
mem[1799] = 8'h90;
mem[1800] = 8'h03;
mem[1801] = 8'h4c;
mem[1802] = 8'h09;
mem[1803] = 8'h07;
mem[1804] = 8'h30;
mem[1805] = 8'h02;
mem[1806] = 8'h10;
mem[1807] = 8'h03;
mem[1808] = 8'h4c;
mem[1809] = 8'h10;
mem[1810] = 8'h07;
mem[1811] = 8'h50;
mem[1812] = 8'h02;
mem[1813] = 8'h70;
mem[1814] = 8'h03;
mem[1815] = 8'h4c;
mem[1816] = 8'h17;
mem[1817] = 8'h07;
mem[1818] = 8'ha9;
mem[1819] = 8'hfd;
mem[1820] = 8'h48;
mem[1821] = 8'h28;
mem[1822] = 8'hf0;
mem[1823] = 8'h02;
mem[1824] = 8'hd0;
mem[1825] = 8'h03;
mem[1826] = 8'h4c;
mem[1827] = 8'h22;
mem[1828] = 8'h07;
mem[1829] = 8'h90;
mem[1830] = 8'h02;
mem[1831] = 8'hb0;
mem[1832] = 8'h03;
mem[1833] = 8'h4c;
mem[1834] = 8'h29;
mem[1835] = 8'h07;
mem[1836] = 8'h10;
mem[1837] = 8'h02;
mem[1838] = 8'h30;
mem[1839] = 8'h03;
mem[1840] = 8'h4c;
mem[1841] = 8'h30;
mem[1842] = 8'h07;
mem[1843] = 8'h50;
mem[1844] = 8'h02;
mem[1845] = 8'h70;
mem[1846] = 8'h03;
mem[1847] = 8'h4c;
mem[1848] = 8'h37;
mem[1849] = 8'h07;
mem[1850] = 8'ha9;
mem[1851] = 8'hfe;
mem[1852] = 8'h48;
mem[1853] = 8'h28;
mem[1854] = 8'hd0;
mem[1855] = 8'h02;
mem[1856] = 8'hf0;
mem[1857] = 8'h03;
mem[1858] = 8'h4c;
mem[1859] = 8'h42;
mem[1860] = 8'h07;
mem[1861] = 8'hb0;
mem[1862] = 8'h02;
mem[1863] = 8'h90;
mem[1864] = 8'h03;
mem[1865] = 8'h4c;
mem[1866] = 8'h49;
mem[1867] = 8'h07;
mem[1868] = 8'h10;
mem[1869] = 8'h02;
mem[1870] = 8'h30;
mem[1871] = 8'h03;
mem[1872] = 8'h4c;
mem[1873] = 8'h50;
mem[1874] = 8'h07;
mem[1875] = 8'h50;
mem[1876] = 8'h02;
mem[1877] = 8'h70;
mem[1878] = 8'h03;
mem[1879] = 8'h4c;
mem[1880] = 8'h57;
mem[1881] = 8'h07;
mem[1882] = 8'ha9;
mem[1883] = 8'h7f;
mem[1884] = 8'h48;
mem[1885] = 8'h28;
mem[1886] = 8'hd0;
mem[1887] = 8'h02;
mem[1888] = 8'hf0;
mem[1889] = 8'h03;
mem[1890] = 8'h4c;
mem[1891] = 8'h62;
mem[1892] = 8'h07;
mem[1893] = 8'h90;
mem[1894] = 8'h02;
mem[1895] = 8'hb0;
mem[1896] = 8'h03;
mem[1897] = 8'h4c;
mem[1898] = 8'h69;
mem[1899] = 8'h07;
mem[1900] = 8'h30;
mem[1901] = 8'h02;
mem[1902] = 8'h10;
mem[1903] = 8'h03;
mem[1904] = 8'h4c;
mem[1905] = 8'h70;
mem[1906] = 8'h07;
mem[1907] = 8'h50;
mem[1908] = 8'h02;
mem[1909] = 8'h70;
mem[1910] = 8'h03;
mem[1911] = 8'h4c;
mem[1912] = 8'h77;
mem[1913] = 8'h07;
mem[1914] = 8'ha9;
mem[1915] = 8'hbf;
mem[1916] = 8'h48;
mem[1917] = 8'h28;
mem[1918] = 8'hd0;
mem[1919] = 8'h02;
mem[1920] = 8'hf0;
mem[1921] = 8'h03;
mem[1922] = 8'h4c;
mem[1923] = 8'h82;
mem[1924] = 8'h07;
mem[1925] = 8'h90;
mem[1926] = 8'h02;
mem[1927] = 8'hb0;
mem[1928] = 8'h03;
mem[1929] = 8'h4c;
mem[1930] = 8'h89;
mem[1931] = 8'h07;
mem[1932] = 8'h10;
mem[1933] = 8'h02;
mem[1934] = 8'h30;
mem[1935] = 8'h03;
mem[1936] = 8'h4c;
mem[1937] = 8'h90;
mem[1938] = 8'h07;
mem[1939] = 8'h70;
mem[1940] = 8'h02;
mem[1941] = 8'h50;
mem[1942] = 8'h03;
mem[1943] = 8'h4c;
mem[1944] = 8'h97;
mem[1945] = 8'h07;
mem[1946] = 8'had;
mem[1947] = 8'h00;
mem[1948] = 8'h02;
mem[1949] = 8'hc9;
mem[1950] = 8'h04;
mem[1951] = 8'hd0;
mem[1952] = 8'hfe;
mem[1953] = 8'ha9;
mem[1954] = 8'h05;
mem[1955] = 8'h8d;
mem[1956] = 8'h00;
mem[1957] = 8'h02;
mem[1958] = 8'ha2;
mem[1959] = 8'h55;
mem[1960] = 8'ha0;
mem[1961] = 8'haa;
mem[1962] = 8'ha9;
mem[1963] = 8'hff;
mem[1964] = 8'h48;
mem[1965] = 8'ha9;
mem[1966] = 8'h01;
mem[1967] = 8'h28;
mem[1968] = 8'h48;
mem[1969] = 8'h08;
mem[1970] = 8'hc9;
mem[1971] = 8'h01;
mem[1972] = 8'hd0;
mem[1973] = 8'hfe;
mem[1974] = 8'h68;
mem[1975] = 8'h48;
mem[1976] = 8'h09;
mem[1977] = 8'h08;
mem[1978] = 8'hc9;
mem[1979] = 8'hff;
mem[1980] = 8'hd0;
mem[1981] = 8'hfe;
mem[1982] = 8'h28;
mem[1983] = 8'ha9;
mem[1984] = 8'h00;
mem[1985] = 8'h48;
mem[1986] = 8'ha9;
mem[1987] = 8'h00;
mem[1988] = 8'h28;
mem[1989] = 8'h48;
mem[1990] = 8'h08;
mem[1991] = 8'hc9;
mem[1992] = 8'h00;
mem[1993] = 8'hd0;
mem[1994] = 8'hfe;
mem[1995] = 8'h68;
mem[1996] = 8'h48;
mem[1997] = 8'h09;
mem[1998] = 8'h08;
mem[1999] = 8'hc9;
mem[2000] = 8'h38;
mem[2001] = 8'hd0;
mem[2002] = 8'hfe;
mem[2003] = 8'h28;
mem[2004] = 8'ha9;
mem[2005] = 8'hff;
mem[2006] = 8'h48;
mem[2007] = 8'ha9;
mem[2008] = 8'hff;
mem[2009] = 8'h28;
mem[2010] = 8'h48;
mem[2011] = 8'h08;
mem[2012] = 8'hc9;
mem[2013] = 8'hff;
mem[2014] = 8'hd0;
mem[2015] = 8'hfe;
mem[2016] = 8'h68;
mem[2017] = 8'h48;
mem[2018] = 8'h09;
mem[2019] = 8'h08;
mem[2020] = 8'hc9;
mem[2021] = 8'hff;
mem[2022] = 8'hd0;
mem[2023] = 8'hfe;
mem[2024] = 8'h28;
mem[2025] = 8'ha9;
mem[2026] = 8'h00;
mem[2027] = 8'h48;
mem[2028] = 8'ha9;
mem[2029] = 8'h01;
mem[2030] = 8'h28;
mem[2031] = 8'h48;
mem[2032] = 8'h08;
mem[2033] = 8'hc9;
mem[2034] = 8'h01;
mem[2035] = 8'hd0;
mem[2036] = 8'hfe;
mem[2037] = 8'h68;
mem[2038] = 8'h48;
mem[2039] = 8'h09;
mem[2040] = 8'h08;
mem[2041] = 8'hc9;
mem[2042] = 8'h38;
mem[2043] = 8'hd0;
mem[2044] = 8'hfe;
mem[2045] = 8'h28;
mem[2046] = 8'ha9;
mem[2047] = 8'hff;
mem[2048] = 8'h48;
mem[2049] = 8'ha9;
mem[2050] = 8'h00;
mem[2051] = 8'h28;
mem[2052] = 8'h48;
mem[2053] = 8'h08;
mem[2054] = 8'hc9;
mem[2055] = 8'h00;
mem[2056] = 8'hd0;
mem[2057] = 8'hfe;
mem[2058] = 8'h68;
mem[2059] = 8'h48;
mem[2060] = 8'h09;
mem[2061] = 8'h08;
mem[2062] = 8'hc9;
mem[2063] = 8'hff;
mem[2064] = 8'hd0;
mem[2065] = 8'hfe;
mem[2066] = 8'h28;
mem[2067] = 8'ha9;
mem[2068] = 8'h00;
mem[2069] = 8'h48;
mem[2070] = 8'ha9;
mem[2071] = 8'hff;
mem[2072] = 8'h28;
mem[2073] = 8'h48;
mem[2074] = 8'h08;
mem[2075] = 8'hc9;
mem[2076] = 8'hff;
mem[2077] = 8'hd0;
mem[2078] = 8'hfe;
mem[2079] = 8'h68;
mem[2080] = 8'h48;
mem[2081] = 8'h09;
mem[2082] = 8'h08;
mem[2083] = 8'hc9;
mem[2084] = 8'h38;
mem[2085] = 8'hd0;
mem[2086] = 8'hfe;
mem[2087] = 8'h28;
mem[2088] = 8'ha9;
mem[2089] = 8'hff;
mem[2090] = 8'h48;
mem[2091] = 8'ha9;
mem[2092] = 8'h00;
mem[2093] = 8'h28;
mem[2094] = 8'h68;
mem[2095] = 8'h08;
mem[2096] = 8'hc9;
mem[2097] = 8'hff;
mem[2098] = 8'hd0;
mem[2099] = 8'hfe;
mem[2100] = 8'h68;
mem[2101] = 8'h48;
mem[2102] = 8'h09;
mem[2103] = 8'h08;
mem[2104] = 8'hc9;
mem[2105] = 8'hfd;
mem[2106] = 8'hd0;
mem[2107] = 8'hfe;
mem[2108] = 8'h28;
mem[2109] = 8'ha9;
mem[2110] = 8'h00;
mem[2111] = 8'h48;
mem[2112] = 8'ha9;
mem[2113] = 8'hff;
mem[2114] = 8'h28;
mem[2115] = 8'h68;
mem[2116] = 8'h08;
mem[2117] = 8'hc9;
mem[2118] = 8'h00;
mem[2119] = 8'hd0;
mem[2120] = 8'hfe;
mem[2121] = 8'h68;
mem[2122] = 8'h48;
mem[2123] = 8'h09;
mem[2124] = 8'h08;
mem[2125] = 8'hc9;
mem[2126] = 8'h3a;
mem[2127] = 8'hd0;
mem[2128] = 8'hfe;
mem[2129] = 8'h28;
mem[2130] = 8'ha9;
mem[2131] = 8'hff;
mem[2132] = 8'h48;
mem[2133] = 8'ha9;
mem[2134] = 8'hfe;
mem[2135] = 8'h28;
mem[2136] = 8'h68;
mem[2137] = 8'h08;
mem[2138] = 8'hc9;
mem[2139] = 8'h01;
mem[2140] = 8'hd0;
mem[2141] = 8'hfe;
mem[2142] = 8'h68;
mem[2143] = 8'h48;
mem[2144] = 8'h09;
mem[2145] = 8'h08;
mem[2146] = 8'hc9;
mem[2147] = 8'h7d;
mem[2148] = 8'hd0;
mem[2149] = 8'hfe;
mem[2150] = 8'h28;
mem[2151] = 8'ha9;
mem[2152] = 8'h00;
mem[2153] = 8'h48;
mem[2154] = 8'ha9;
mem[2155] = 8'h00;
mem[2156] = 8'h28;
mem[2157] = 8'h68;
mem[2158] = 8'h08;
mem[2159] = 8'hc9;
mem[2160] = 8'hff;
mem[2161] = 8'hd0;
mem[2162] = 8'hfe;
mem[2163] = 8'h68;
mem[2164] = 8'h48;
mem[2165] = 8'h09;
mem[2166] = 8'h08;
mem[2167] = 8'hc9;
mem[2168] = 8'hb8;
mem[2169] = 8'hd0;
mem[2170] = 8'hfe;
mem[2171] = 8'h28;
mem[2172] = 8'ha9;
mem[2173] = 8'hff;
mem[2174] = 8'h48;
mem[2175] = 8'ha9;
mem[2176] = 8'hff;
mem[2177] = 8'h28;
mem[2178] = 8'h68;
mem[2179] = 8'h08;
mem[2180] = 8'hc9;
mem[2181] = 8'h00;
mem[2182] = 8'hd0;
mem[2183] = 8'hfe;
mem[2184] = 8'h68;
mem[2185] = 8'h48;
mem[2186] = 8'h09;
mem[2187] = 8'h08;
mem[2188] = 8'hc9;
mem[2189] = 8'h7f;
mem[2190] = 8'hd0;
mem[2191] = 8'hfe;
mem[2192] = 8'h28;
mem[2193] = 8'ha9;
mem[2194] = 8'h00;
mem[2195] = 8'h48;
mem[2196] = 8'ha9;
mem[2197] = 8'hfe;
mem[2198] = 8'h28;
mem[2199] = 8'h68;
mem[2200] = 8'h08;
mem[2201] = 8'hc9;
mem[2202] = 8'h01;
mem[2203] = 8'hd0;
mem[2204] = 8'hfe;
mem[2205] = 8'h68;
mem[2206] = 8'h48;
mem[2207] = 8'h09;
mem[2208] = 8'h08;
mem[2209] = 8'hc9;
mem[2210] = 8'h38;
mem[2211] = 8'hd0;
mem[2212] = 8'hfe;
mem[2213] = 8'h28;
mem[2214] = 8'he0;
mem[2215] = 8'h55;
mem[2216] = 8'hd0;
mem[2217] = 8'hfe;
mem[2218] = 8'hc0;
mem[2219] = 8'haa;
mem[2220] = 8'hd0;
mem[2221] = 8'hfe;
mem[2222] = 8'had;
mem[2223] = 8'h00;
mem[2224] = 8'h02;
mem[2225] = 8'hc9;
mem[2226] = 8'h05;
mem[2227] = 8'hd0;
mem[2228] = 8'hfe;
mem[2229] = 8'ha9;
mem[2230] = 8'h06;
mem[2231] = 8'h8d;
mem[2232] = 8'h00;
mem[2233] = 8'h02;
mem[2234] = 8'ha9;
mem[2235] = 8'h00;
mem[2236] = 8'h48;
mem[2237] = 8'ha9;
mem[2238] = 8'h3c;
mem[2239] = 8'h28;
mem[2240] = 8'h49;
mem[2241] = 8'hc3;
mem[2242] = 8'h08;
mem[2243] = 8'hc9;
mem[2244] = 8'hff;
mem[2245] = 8'hd0;
mem[2246] = 8'hfe;
mem[2247] = 8'h68;
mem[2248] = 8'h48;
mem[2249] = 8'h09;
mem[2250] = 8'h08;
mem[2251] = 8'hc9;
mem[2252] = 8'hb8;
mem[2253] = 8'hd0;
mem[2254] = 8'hfe;
mem[2255] = 8'h28;
mem[2256] = 8'ha9;
mem[2257] = 8'h00;
mem[2258] = 8'h48;
mem[2259] = 8'ha9;
mem[2260] = 8'hc3;
mem[2261] = 8'h28;
mem[2262] = 8'h49;
mem[2263] = 8'hc3;
mem[2264] = 8'h08;
mem[2265] = 8'hc9;
mem[2266] = 8'h00;
mem[2267] = 8'hd0;
mem[2268] = 8'hfe;
mem[2269] = 8'h68;
mem[2270] = 8'h48;
mem[2271] = 8'h09;
mem[2272] = 8'h08;
mem[2273] = 8'hc9;
mem[2274] = 8'h3a;
mem[2275] = 8'hd0;
mem[2276] = 8'hfe;
mem[2277] = 8'h28;
mem[2278] = 8'had;
mem[2279] = 8'h00;
mem[2280] = 8'h02;
mem[2281] = 8'hc9;
mem[2282] = 8'h06;
mem[2283] = 8'hd0;
mem[2284] = 8'hfe;
mem[2285] = 8'ha9;
mem[2286] = 8'h07;
mem[2287] = 8'h8d;
mem[2288] = 8'h00;
mem[2289] = 8'h02;
mem[2290] = 8'ha2;
mem[2291] = 8'h24;
mem[2292] = 8'ha0;
mem[2293] = 8'h42;
mem[2294] = 8'ha9;
mem[2295] = 8'h00;
mem[2296] = 8'h48;
mem[2297] = 8'ha9;
mem[2298] = 8'h18;
mem[2299] = 8'h28;
mem[2300] = 8'hea;
mem[2301] = 8'h08;
mem[2302] = 8'hc9;
mem[2303] = 8'h18;
mem[2304] = 8'hd0;
mem[2305] = 8'hfe;
mem[2306] = 8'h68;
mem[2307] = 8'h48;
mem[2308] = 8'h09;
mem[2309] = 8'h08;
mem[2310] = 8'hc9;
mem[2311] = 8'h38;
mem[2312] = 8'hd0;
mem[2313] = 8'hfe;
mem[2314] = 8'h28;
mem[2315] = 8'he0;
mem[2316] = 8'h24;
mem[2317] = 8'hd0;
mem[2318] = 8'hfe;
mem[2319] = 8'hc0;
mem[2320] = 8'h42;
mem[2321] = 8'hd0;
mem[2322] = 8'hfe;
mem[2323] = 8'ha2;
mem[2324] = 8'hdb;
mem[2325] = 8'ha0;
mem[2326] = 8'hbd;
mem[2327] = 8'ha9;
mem[2328] = 8'hff;
mem[2329] = 8'h48;
mem[2330] = 8'ha9;
mem[2331] = 8'he7;
mem[2332] = 8'h28;
mem[2333] = 8'hea;
mem[2334] = 8'h08;
mem[2335] = 8'hc9;
mem[2336] = 8'he7;
mem[2337] = 8'hd0;
mem[2338] = 8'hfe;
mem[2339] = 8'h68;
mem[2340] = 8'h48;
mem[2341] = 8'h09;
mem[2342] = 8'h08;
mem[2343] = 8'hc9;
mem[2344] = 8'hff;
mem[2345] = 8'hd0;
mem[2346] = 8'hfe;
mem[2347] = 8'h28;
mem[2348] = 8'he0;
mem[2349] = 8'hdb;
mem[2350] = 8'hd0;
mem[2351] = 8'hfe;
mem[2352] = 8'hc0;
mem[2353] = 8'hbd;
mem[2354] = 8'hd0;
mem[2355] = 8'hfe;
mem[2356] = 8'had;
mem[2357] = 8'h00;
mem[2358] = 8'h02;
mem[2359] = 8'hc9;
mem[2360] = 8'h07;
mem[2361] = 8'hd0;
mem[2362] = 8'hfe;
mem[2363] = 8'ha9;
mem[2364] = 8'h08;
mem[2365] = 8'h8d;
mem[2366] = 8'h00;
mem[2367] = 8'h02;
mem[2368] = 8'ha9;
mem[2369] = 8'h00;
mem[2370] = 8'h48;
mem[2371] = 8'h28;
mem[2372] = 8'ha9;
mem[2373] = 8'h46;
mem[2374] = 8'ha2;
mem[2375] = 8'h41;
mem[2376] = 8'ha0;
mem[2377] = 8'h52;
mem[2378] = 8'h4c;
mem[2379] = 8'he4;
mem[2380] = 8'h37;
mem[2381] = 8'hea;
mem[2382] = 8'hea;
mem[2383] = 8'hd0;
mem[2384] = 8'hfe;
mem[2385] = 8'he8;
mem[2386] = 8'he8;
mem[2387] = 8'hf0;
mem[2388] = 8'hfe;
mem[2389] = 8'h10;
mem[2390] = 8'hfe;
mem[2391] = 8'h90;
mem[2392] = 8'hfe;
mem[2393] = 8'h50;
mem[2394] = 8'hfe;
mem[2395] = 8'hc9;
mem[2396] = 8'hec;
mem[2397] = 8'hd0;
mem[2398] = 8'hfe;
mem[2399] = 8'he0;
mem[2400] = 8'h42;
mem[2401] = 8'hd0;
mem[2402] = 8'hfe;
mem[2403] = 8'hc0;
mem[2404] = 8'h4f;
mem[2405] = 8'hd0;
mem[2406] = 8'hfe;
mem[2407] = 8'hca;
mem[2408] = 8'hc8;
mem[2409] = 8'hc8;
mem[2410] = 8'hc8;
mem[2411] = 8'h49;
mem[2412] = 8'haa;
mem[2413] = 8'h4c;
mem[2414] = 8'h76;
mem[2415] = 8'h09;
mem[2416] = 8'hea;
mem[2417] = 8'hea;
mem[2418] = 8'hd0;
mem[2419] = 8'hfe;
mem[2420] = 8'he8;
mem[2421] = 8'he8;
mem[2422] = 8'hf0;
mem[2423] = 8'hfe;
mem[2424] = 8'h30;
mem[2425] = 8'hfe;
mem[2426] = 8'h90;
mem[2427] = 8'hfe;
mem[2428] = 8'h50;
mem[2429] = 8'hfe;
mem[2430] = 8'hc9;
mem[2431] = 8'h46;
mem[2432] = 8'hd0;
mem[2433] = 8'hfe;
mem[2434] = 8'he0;
mem[2435] = 8'h41;
mem[2436] = 8'hd0;
mem[2437] = 8'hfe;
mem[2438] = 8'hc0;
mem[2439] = 8'h52;
mem[2440] = 8'hd0;
mem[2441] = 8'hfe;
mem[2442] = 8'had;
mem[2443] = 8'h00;
mem[2444] = 8'h02;
mem[2445] = 8'hc9;
mem[2446] = 8'h08;
mem[2447] = 8'hd0;
mem[2448] = 8'hfe;
mem[2449] = 8'ha9;
mem[2450] = 8'h09;
mem[2451] = 8'h8d;
mem[2452] = 8'h00;
mem[2453] = 8'h02;
mem[2454] = 8'ha9;
mem[2455] = 8'h00;
mem[2456] = 8'h48;
mem[2457] = 8'h28;
mem[2458] = 8'ha9;
mem[2459] = 8'h49;
mem[2460] = 8'ha2;
mem[2461] = 8'h4e;
mem[2462] = 8'ha0;
mem[2463] = 8'h44;
mem[2464] = 8'h6c;
mem[2465] = 8'h12;
mem[2466] = 8'h38;
mem[2467] = 8'hea;
mem[2468] = 8'hd0;
mem[2469] = 8'hfe;
mem[2470] = 8'h88;
mem[2471] = 8'h88;
mem[2472] = 8'h08;
mem[2473] = 8'h88;
mem[2474] = 8'h88;
mem[2475] = 8'h88;
mem[2476] = 8'h28;
mem[2477] = 8'hf0;
mem[2478] = 8'hfe;
mem[2479] = 8'h10;
mem[2480] = 8'hfe;
mem[2481] = 8'h90;
mem[2482] = 8'hfe;
mem[2483] = 8'h50;
mem[2484] = 8'hfe;
mem[2485] = 8'hc9;
mem[2486] = 8'he3;
mem[2487] = 8'hd0;
mem[2488] = 8'hfe;
mem[2489] = 8'he0;
mem[2490] = 8'h4f;
mem[2491] = 8'hd0;
mem[2492] = 8'hfe;
mem[2493] = 8'hc0;
mem[2494] = 8'h3e;
mem[2495] = 8'hd0;
mem[2496] = 8'hfe;
mem[2497] = 8'hba;
mem[2498] = 8'he0;
mem[2499] = 8'hff;
mem[2500] = 8'hd0;
mem[2501] = 8'hfe;
mem[2502] = 8'had;
mem[2503] = 8'h00;
mem[2504] = 8'h02;
mem[2505] = 8'hc9;
mem[2506] = 8'h09;
mem[2507] = 8'hd0;
mem[2508] = 8'hfe;
mem[2509] = 8'ha9;
mem[2510] = 8'h0a;
mem[2511] = 8'h8d;
mem[2512] = 8'h00;
mem[2513] = 8'h02;
mem[2514] = 8'ha9;
mem[2515] = 8'h00;
mem[2516] = 8'h48;
mem[2517] = 8'h28;
mem[2518] = 8'ha9;
mem[2519] = 8'h4a;
mem[2520] = 8'ha2;
mem[2521] = 8'h53;
mem[2522] = 8'ha0;
mem[2523] = 8'h52;
mem[2524] = 8'h20;
mem[2525] = 8'h4e;
mem[2526] = 8'h38;
mem[2527] = 8'h08;
mem[2528] = 8'h88;
mem[2529] = 8'h88;
mem[2530] = 8'h88;
mem[2531] = 8'h28;
mem[2532] = 8'hf0;
mem[2533] = 8'hfe;
mem[2534] = 8'h10;
mem[2535] = 8'hfe;
mem[2536] = 8'h90;
mem[2537] = 8'hfe;
mem[2538] = 8'h50;
mem[2539] = 8'hfe;
mem[2540] = 8'hc9;
mem[2541] = 8'he0;
mem[2542] = 8'hd0;
mem[2543] = 8'hfe;
mem[2544] = 8'he0;
mem[2545] = 8'h54;
mem[2546] = 8'hd0;
mem[2547] = 8'hfe;
mem[2548] = 8'hc0;
mem[2549] = 8'h4c;
mem[2550] = 8'hd0;
mem[2551] = 8'hfe;
mem[2552] = 8'hba;
mem[2553] = 8'he0;
mem[2554] = 8'hff;
mem[2555] = 8'hd0;
mem[2556] = 8'hfe;
mem[2557] = 8'had;
mem[2558] = 8'h00;
mem[2559] = 8'h02;
mem[2560] = 8'hc9;
mem[2561] = 8'h0a;
mem[2562] = 8'hd0;
mem[2563] = 8'hfe;
mem[2564] = 8'ha9;
mem[2565] = 8'h0b;
mem[2566] = 8'h8d;
mem[2567] = 8'h00;
mem[2568] = 8'h02;
mem[2569] = 8'ha9;
mem[2570] = 8'h00;
mem[2571] = 8'h48;
mem[2572] = 8'h28;
mem[2573] = 8'ha9;
mem[2574] = 8'h42;
mem[2575] = 8'ha2;
mem[2576] = 8'h52;
mem[2577] = 8'ha0;
mem[2578] = 8'h4b;
mem[2579] = 8'h00;
mem[2580] = 8'h88;
mem[2581] = 8'h08;
mem[2582] = 8'h88;
mem[2583] = 8'h88;
mem[2584] = 8'h88;
mem[2585] = 8'hc9;
mem[2586] = 8'he8;
mem[2587] = 8'hd0;
mem[2588] = 8'hfe;
mem[2589] = 8'he0;
mem[2590] = 8'h53;
mem[2591] = 8'hd0;
mem[2592] = 8'hfe;
mem[2593] = 8'hc0;
mem[2594] = 8'h45;
mem[2595] = 8'hd0;
mem[2596] = 8'hfe;
mem[2597] = 8'h68;
mem[2598] = 8'h09;
mem[2599] = 8'h08;
mem[2600] = 8'hc9;
mem[2601] = 8'h38;
mem[2602] = 8'hd0;
mem[2603] = 8'hfe;
mem[2604] = 8'hba;
mem[2605] = 8'he0;
mem[2606] = 8'hff;
mem[2607] = 8'hd0;
mem[2608] = 8'hfe;
mem[2609] = 8'had;
mem[2610] = 8'h00;
mem[2611] = 8'h02;
mem[2612] = 8'hc9;
mem[2613] = 8'h0b;
mem[2614] = 8'hd0;
mem[2615] = 8'hfe;
mem[2616] = 8'ha9;
mem[2617] = 8'h0c;
mem[2618] = 8'h8d;
mem[2619] = 8'h00;
mem[2620] = 8'h02;
mem[2621] = 8'ha9;
mem[2622] = 8'hff;
mem[2623] = 8'h48;
mem[2624] = 8'h28;
mem[2625] = 8'h18;
mem[2626] = 8'h08;
mem[2627] = 8'h68;
mem[2628] = 8'h48;
mem[2629] = 8'h09;
mem[2630] = 8'h08;
mem[2631] = 8'hc9;
mem[2632] = 8'hfe;
mem[2633] = 8'hd0;
mem[2634] = 8'hfe;
mem[2635] = 8'h28;
mem[2636] = 8'h38;
mem[2637] = 8'h08;
mem[2638] = 8'h68;
mem[2639] = 8'h48;
mem[2640] = 8'h09;
mem[2641] = 8'h08;
mem[2642] = 8'hc9;
mem[2643] = 8'hff;
mem[2644] = 8'hd0;
mem[2645] = 8'hfe;
mem[2646] = 8'h28;
mem[2647] = 8'h58;
mem[2648] = 8'h08;
mem[2649] = 8'h68;
mem[2650] = 8'h48;
mem[2651] = 8'h09;
mem[2652] = 8'h08;
mem[2653] = 8'hc9;
mem[2654] = 8'hfb;
mem[2655] = 8'hd0;
mem[2656] = 8'hfe;
mem[2657] = 8'h28;
mem[2658] = 8'h78;
mem[2659] = 8'h08;
mem[2660] = 8'h68;
mem[2661] = 8'h48;
mem[2662] = 8'h09;
mem[2663] = 8'h08;
mem[2664] = 8'hc9;
mem[2665] = 8'hff;
mem[2666] = 8'hd0;
mem[2667] = 8'hfe;
mem[2668] = 8'h28;
mem[2669] = 8'hd8;
mem[2670] = 8'h08;
mem[2671] = 8'h68;
mem[2672] = 8'h48;
mem[2673] = 8'h09;
mem[2674] = 8'h08;
mem[2675] = 8'hc9;
mem[2676] = 8'hff;
mem[2677] = 8'hd0;
mem[2678] = 8'hfe;
mem[2679] = 8'h28;
mem[2680] = 8'hf8;
mem[2681] = 8'h08;
mem[2682] = 8'h68;
mem[2683] = 8'h48;
mem[2684] = 8'h09;
mem[2685] = 8'h08;
mem[2686] = 8'hc9;
mem[2687] = 8'hff;
mem[2688] = 8'hd0;
mem[2689] = 8'hfe;
mem[2690] = 8'h28;
mem[2691] = 8'hb8;
mem[2692] = 8'h08;
mem[2693] = 8'h68;
mem[2694] = 8'h48;
mem[2695] = 8'h09;
mem[2696] = 8'h08;
mem[2697] = 8'hc9;
mem[2698] = 8'hbf;
mem[2699] = 8'hd0;
mem[2700] = 8'hfe;
mem[2701] = 8'h28;
mem[2702] = 8'ha9;
mem[2703] = 8'h00;
mem[2704] = 8'h48;
mem[2705] = 8'h28;
mem[2706] = 8'h08;
mem[2707] = 8'h68;
mem[2708] = 8'h48;
mem[2709] = 8'h09;
mem[2710] = 8'h08;
mem[2711] = 8'hc9;
mem[2712] = 8'h38;
mem[2713] = 8'hd0;
mem[2714] = 8'hfe;
mem[2715] = 8'h28;
mem[2716] = 8'h38;
mem[2717] = 8'h08;
mem[2718] = 8'h68;
mem[2719] = 8'h48;
mem[2720] = 8'h09;
mem[2721] = 8'h08;
mem[2722] = 8'hc9;
mem[2723] = 8'h39;
mem[2724] = 8'hd0;
mem[2725] = 8'hfe;
mem[2726] = 8'h28;
mem[2727] = 8'h18;
mem[2728] = 8'h08;
mem[2729] = 8'h68;
mem[2730] = 8'h48;
mem[2731] = 8'h09;
mem[2732] = 8'h08;
mem[2733] = 8'hc9;
mem[2734] = 8'h38;
mem[2735] = 8'hd0;
mem[2736] = 8'hfe;
mem[2737] = 8'h28;
mem[2738] = 8'h78;
mem[2739] = 8'h08;
mem[2740] = 8'h68;
mem[2741] = 8'h48;
mem[2742] = 8'h09;
mem[2743] = 8'h08;
mem[2744] = 8'hc9;
mem[2745] = 8'h3c;
mem[2746] = 8'hd0;
mem[2747] = 8'hfe;
mem[2748] = 8'h28;
mem[2749] = 8'h58;
mem[2750] = 8'h08;
mem[2751] = 8'h68;
mem[2752] = 8'h48;
mem[2753] = 8'h09;
mem[2754] = 8'h08;
mem[2755] = 8'hc9;
mem[2756] = 8'h38;
mem[2757] = 8'hd0;
mem[2758] = 8'hfe;
mem[2759] = 8'h28;
mem[2760] = 8'hf8;
mem[2761] = 8'h08;
mem[2762] = 8'h68;
mem[2763] = 8'h48;
mem[2764] = 8'h09;
mem[2765] = 8'h08;
mem[2766] = 8'hc9;
mem[2767] = 8'h38;
mem[2768] = 8'hd0;
mem[2769] = 8'hfe;
mem[2770] = 8'h28;
mem[2771] = 8'hd8;
mem[2772] = 8'h08;
mem[2773] = 8'h68;
mem[2774] = 8'h48;
mem[2775] = 8'h09;
mem[2776] = 8'h08;
mem[2777] = 8'hc9;
mem[2778] = 8'h38;
mem[2779] = 8'hd0;
mem[2780] = 8'hfe;
mem[2781] = 8'h28;
mem[2782] = 8'ha9;
mem[2783] = 8'h40;
mem[2784] = 8'h48;
mem[2785] = 8'h28;
mem[2786] = 8'h08;
mem[2787] = 8'h68;
mem[2788] = 8'h48;
mem[2789] = 8'h09;
mem[2790] = 8'h08;
mem[2791] = 8'hc9;
mem[2792] = 8'h78;
mem[2793] = 8'hd0;
mem[2794] = 8'hfe;
mem[2795] = 8'h28;
mem[2796] = 8'hb8;
mem[2797] = 8'h08;
mem[2798] = 8'h68;
mem[2799] = 8'h48;
mem[2800] = 8'h09;
mem[2801] = 8'h08;
mem[2802] = 8'hc9;
mem[2803] = 8'h38;
mem[2804] = 8'hd0;
mem[2805] = 8'hfe;
mem[2806] = 8'h28;
mem[2807] = 8'had;
mem[2808] = 8'h00;
mem[2809] = 8'h02;
mem[2810] = 8'hc9;
mem[2811] = 8'h0c;
mem[2812] = 8'hd0;
mem[2813] = 8'hfe;
mem[2814] = 8'ha9;
mem[2815] = 8'h0d;
mem[2816] = 8'h8d;
mem[2817] = 8'h00;
mem[2818] = 8'h02;
mem[2819] = 8'ha2;
mem[2820] = 8'hfe;
mem[2821] = 8'ha9;
mem[2822] = 8'hff;
mem[2823] = 8'h48;
mem[2824] = 8'h28;
mem[2825] = 8'he8;
mem[2826] = 8'h08;
mem[2827] = 8'he0;
mem[2828] = 8'hff;
mem[2829] = 8'hd0;
mem[2830] = 8'hfe;
mem[2831] = 8'h68;
mem[2832] = 8'h48;
mem[2833] = 8'h09;
mem[2834] = 8'h08;
mem[2835] = 8'hc9;
mem[2836] = 8'hfd;
mem[2837] = 8'hd0;
mem[2838] = 8'hfe;
mem[2839] = 8'h28;
mem[2840] = 8'he8;
mem[2841] = 8'h08;
mem[2842] = 8'he0;
mem[2843] = 8'h00;
mem[2844] = 8'hd0;
mem[2845] = 8'hfe;
mem[2846] = 8'h68;
mem[2847] = 8'h48;
mem[2848] = 8'h09;
mem[2849] = 8'h08;
mem[2850] = 8'hc9;
mem[2851] = 8'h7f;
mem[2852] = 8'hd0;
mem[2853] = 8'hfe;
mem[2854] = 8'h28;
mem[2855] = 8'he8;
mem[2856] = 8'h08;
mem[2857] = 8'he0;
mem[2858] = 8'h01;
mem[2859] = 8'hd0;
mem[2860] = 8'hfe;
mem[2861] = 8'h68;
mem[2862] = 8'h48;
mem[2863] = 8'h09;
mem[2864] = 8'h08;
mem[2865] = 8'hc9;
mem[2866] = 8'h7d;
mem[2867] = 8'hd0;
mem[2868] = 8'hfe;
mem[2869] = 8'h28;
mem[2870] = 8'hca;
mem[2871] = 8'h08;
mem[2872] = 8'he0;
mem[2873] = 8'h00;
mem[2874] = 8'hd0;
mem[2875] = 8'hfe;
mem[2876] = 8'h68;
mem[2877] = 8'h48;
mem[2878] = 8'h09;
mem[2879] = 8'h08;
mem[2880] = 8'hc9;
mem[2881] = 8'h7f;
mem[2882] = 8'hd0;
mem[2883] = 8'hfe;
mem[2884] = 8'h28;
mem[2885] = 8'hca;
mem[2886] = 8'h08;
mem[2887] = 8'he0;
mem[2888] = 8'hff;
mem[2889] = 8'hd0;
mem[2890] = 8'hfe;
mem[2891] = 8'h68;
mem[2892] = 8'h48;
mem[2893] = 8'h09;
mem[2894] = 8'h08;
mem[2895] = 8'hc9;
mem[2896] = 8'hfd;
mem[2897] = 8'hd0;
mem[2898] = 8'hfe;
mem[2899] = 8'h28;
mem[2900] = 8'hca;
mem[2901] = 8'ha9;
mem[2902] = 8'h00;
mem[2903] = 8'h48;
mem[2904] = 8'h28;
mem[2905] = 8'he8;
mem[2906] = 8'h08;
mem[2907] = 8'he0;
mem[2908] = 8'hff;
mem[2909] = 8'hd0;
mem[2910] = 8'hfe;
mem[2911] = 8'h68;
mem[2912] = 8'h48;
mem[2913] = 8'h09;
mem[2914] = 8'h08;
mem[2915] = 8'hc9;
mem[2916] = 8'hb8;
mem[2917] = 8'hd0;
mem[2918] = 8'hfe;
mem[2919] = 8'h28;
mem[2920] = 8'he8;
mem[2921] = 8'h08;
mem[2922] = 8'he0;
mem[2923] = 8'h00;
mem[2924] = 8'hd0;
mem[2925] = 8'hfe;
mem[2926] = 8'h68;
mem[2927] = 8'h48;
mem[2928] = 8'h09;
mem[2929] = 8'h08;
mem[2930] = 8'hc9;
mem[2931] = 8'h3a;
mem[2932] = 8'hd0;
mem[2933] = 8'hfe;
mem[2934] = 8'h28;
mem[2935] = 8'he8;
mem[2936] = 8'h08;
mem[2937] = 8'he0;
mem[2938] = 8'h01;
mem[2939] = 8'hd0;
mem[2940] = 8'hfe;
mem[2941] = 8'h68;
mem[2942] = 8'h48;
mem[2943] = 8'h09;
mem[2944] = 8'h08;
mem[2945] = 8'hc9;
mem[2946] = 8'h38;
mem[2947] = 8'hd0;
mem[2948] = 8'hfe;
mem[2949] = 8'h28;
mem[2950] = 8'hca;
mem[2951] = 8'h08;
mem[2952] = 8'he0;
mem[2953] = 8'h00;
mem[2954] = 8'hd0;
mem[2955] = 8'hfe;
mem[2956] = 8'h68;
mem[2957] = 8'h48;
mem[2958] = 8'h09;
mem[2959] = 8'h08;
mem[2960] = 8'hc9;
mem[2961] = 8'h3a;
mem[2962] = 8'hd0;
mem[2963] = 8'hfe;
mem[2964] = 8'h28;
mem[2965] = 8'hca;
mem[2966] = 8'h08;
mem[2967] = 8'he0;
mem[2968] = 8'hff;
mem[2969] = 8'hd0;
mem[2970] = 8'hfe;
mem[2971] = 8'h68;
mem[2972] = 8'h48;
mem[2973] = 8'h09;
mem[2974] = 8'h08;
mem[2975] = 8'hc9;
mem[2976] = 8'hb8;
mem[2977] = 8'hd0;
mem[2978] = 8'hfe;
mem[2979] = 8'h28;
mem[2980] = 8'ha0;
mem[2981] = 8'hfe;
mem[2982] = 8'ha9;
mem[2983] = 8'hff;
mem[2984] = 8'h48;
mem[2985] = 8'h28;
mem[2986] = 8'hc8;
mem[2987] = 8'h08;
mem[2988] = 8'hc0;
mem[2989] = 8'hff;
mem[2990] = 8'hd0;
mem[2991] = 8'hfe;
mem[2992] = 8'h68;
mem[2993] = 8'h48;
mem[2994] = 8'h09;
mem[2995] = 8'h08;
mem[2996] = 8'hc9;
mem[2997] = 8'hfd;
mem[2998] = 8'hd0;
mem[2999] = 8'hfe;
mem[3000] = 8'h28;
mem[3001] = 8'hc8;
mem[3002] = 8'h08;
mem[3003] = 8'hc0;
mem[3004] = 8'h00;
mem[3005] = 8'hd0;
mem[3006] = 8'hfe;
mem[3007] = 8'h68;
mem[3008] = 8'h48;
mem[3009] = 8'h09;
mem[3010] = 8'h08;
mem[3011] = 8'hc9;
mem[3012] = 8'h7f;
mem[3013] = 8'hd0;
mem[3014] = 8'hfe;
mem[3015] = 8'h28;
mem[3016] = 8'hc8;
mem[3017] = 8'h08;
mem[3018] = 8'hc0;
mem[3019] = 8'h01;
mem[3020] = 8'hd0;
mem[3021] = 8'hfe;
mem[3022] = 8'h68;
mem[3023] = 8'h48;
mem[3024] = 8'h09;
mem[3025] = 8'h08;
mem[3026] = 8'hc9;
mem[3027] = 8'h7d;
mem[3028] = 8'hd0;
mem[3029] = 8'hfe;
mem[3030] = 8'h28;
mem[3031] = 8'h88;
mem[3032] = 8'h08;
mem[3033] = 8'hc0;
mem[3034] = 8'h00;
mem[3035] = 8'hd0;
mem[3036] = 8'hfe;
mem[3037] = 8'h68;
mem[3038] = 8'h48;
mem[3039] = 8'h09;
mem[3040] = 8'h08;
mem[3041] = 8'hc9;
mem[3042] = 8'h7f;
mem[3043] = 8'hd0;
mem[3044] = 8'hfe;
mem[3045] = 8'h28;
mem[3046] = 8'h88;
mem[3047] = 8'h08;
mem[3048] = 8'hc0;
mem[3049] = 8'hff;
mem[3050] = 8'hd0;
mem[3051] = 8'hfe;
mem[3052] = 8'h68;
mem[3053] = 8'h48;
mem[3054] = 8'h09;
mem[3055] = 8'h08;
mem[3056] = 8'hc9;
mem[3057] = 8'hfd;
mem[3058] = 8'hd0;
mem[3059] = 8'hfe;
mem[3060] = 8'h28;
mem[3061] = 8'h88;
mem[3062] = 8'ha9;
mem[3063] = 8'h00;
mem[3064] = 8'h48;
mem[3065] = 8'h28;
mem[3066] = 8'hc8;
mem[3067] = 8'h08;
mem[3068] = 8'hc0;
mem[3069] = 8'hff;
mem[3070] = 8'hd0;
mem[3071] = 8'hfe;
mem[3072] = 8'h68;
mem[3073] = 8'h48;
mem[3074] = 8'h09;
mem[3075] = 8'h08;
mem[3076] = 8'hc9;
mem[3077] = 8'hb8;
mem[3078] = 8'hd0;
mem[3079] = 8'hfe;
mem[3080] = 8'h28;
mem[3081] = 8'hc8;
mem[3082] = 8'h08;
mem[3083] = 8'hc0;
mem[3084] = 8'h00;
mem[3085] = 8'hd0;
mem[3086] = 8'hfe;
mem[3087] = 8'h68;
mem[3088] = 8'h48;
mem[3089] = 8'h09;
mem[3090] = 8'h08;
mem[3091] = 8'hc9;
mem[3092] = 8'h3a;
mem[3093] = 8'hd0;
mem[3094] = 8'hfe;
mem[3095] = 8'h28;
mem[3096] = 8'hc8;
mem[3097] = 8'h08;
mem[3098] = 8'hc0;
mem[3099] = 8'h01;
mem[3100] = 8'hd0;
mem[3101] = 8'hfe;
mem[3102] = 8'h68;
mem[3103] = 8'h48;
mem[3104] = 8'h09;
mem[3105] = 8'h08;
mem[3106] = 8'hc9;
mem[3107] = 8'h38;
mem[3108] = 8'hd0;
mem[3109] = 8'hfe;
mem[3110] = 8'h28;
mem[3111] = 8'h88;
mem[3112] = 8'h08;
mem[3113] = 8'hc0;
mem[3114] = 8'h00;
mem[3115] = 8'hd0;
mem[3116] = 8'hfe;
mem[3117] = 8'h68;
mem[3118] = 8'h48;
mem[3119] = 8'h09;
mem[3120] = 8'h08;
mem[3121] = 8'hc9;
mem[3122] = 8'h3a;
mem[3123] = 8'hd0;
mem[3124] = 8'hfe;
mem[3125] = 8'h28;
mem[3126] = 8'h88;
mem[3127] = 8'h08;
mem[3128] = 8'hc0;
mem[3129] = 8'hff;
mem[3130] = 8'hd0;
mem[3131] = 8'hfe;
mem[3132] = 8'h68;
mem[3133] = 8'h48;
mem[3134] = 8'h09;
mem[3135] = 8'h08;
mem[3136] = 8'hc9;
mem[3137] = 8'hb8;
mem[3138] = 8'hd0;
mem[3139] = 8'hfe;
mem[3140] = 8'h28;
mem[3141] = 8'ha2;
mem[3142] = 8'hff;
mem[3143] = 8'ha9;
mem[3144] = 8'hff;
mem[3145] = 8'h48;
mem[3146] = 8'h28;
mem[3147] = 8'h8a;
mem[3148] = 8'h08;
mem[3149] = 8'hc9;
mem[3150] = 8'hff;
mem[3151] = 8'hd0;
mem[3152] = 8'hfe;
mem[3153] = 8'h68;
mem[3154] = 8'h48;
mem[3155] = 8'h09;
mem[3156] = 8'h08;
mem[3157] = 8'hc9;
mem[3158] = 8'hfd;
mem[3159] = 8'hd0;
mem[3160] = 8'hfe;
mem[3161] = 8'h28;
mem[3162] = 8'h08;
mem[3163] = 8'he8;
mem[3164] = 8'h28;
mem[3165] = 8'h8a;
mem[3166] = 8'h08;
mem[3167] = 8'hc9;
mem[3168] = 8'h00;
mem[3169] = 8'hd0;
mem[3170] = 8'hfe;
mem[3171] = 8'h68;
mem[3172] = 8'h48;
mem[3173] = 8'h09;
mem[3174] = 8'h08;
mem[3175] = 8'hc9;
mem[3176] = 8'h7f;
mem[3177] = 8'hd0;
mem[3178] = 8'hfe;
mem[3179] = 8'h28;
mem[3180] = 8'h08;
mem[3181] = 8'he8;
mem[3182] = 8'h28;
mem[3183] = 8'h8a;
mem[3184] = 8'h08;
mem[3185] = 8'hc9;
mem[3186] = 8'h01;
mem[3187] = 8'hd0;
mem[3188] = 8'hfe;
mem[3189] = 8'h68;
mem[3190] = 8'h48;
mem[3191] = 8'h09;
mem[3192] = 8'h08;
mem[3193] = 8'hc9;
mem[3194] = 8'h7d;
mem[3195] = 8'hd0;
mem[3196] = 8'hfe;
mem[3197] = 8'h28;
mem[3198] = 8'ha9;
mem[3199] = 8'h00;
mem[3200] = 8'h48;
mem[3201] = 8'h28;
mem[3202] = 8'h8a;
mem[3203] = 8'h08;
mem[3204] = 8'hc9;
mem[3205] = 8'h01;
mem[3206] = 8'hd0;
mem[3207] = 8'hfe;
mem[3208] = 8'h68;
mem[3209] = 8'h48;
mem[3210] = 8'h09;
mem[3211] = 8'h08;
mem[3212] = 8'hc9;
mem[3213] = 8'h38;
mem[3214] = 8'hd0;
mem[3215] = 8'hfe;
mem[3216] = 8'h28;
mem[3217] = 8'h08;
mem[3218] = 8'hca;
mem[3219] = 8'h28;
mem[3220] = 8'h8a;
mem[3221] = 8'h08;
mem[3222] = 8'hc9;
mem[3223] = 8'h00;
mem[3224] = 8'hd0;
mem[3225] = 8'hfe;
mem[3226] = 8'h68;
mem[3227] = 8'h48;
mem[3228] = 8'h09;
mem[3229] = 8'h08;
mem[3230] = 8'hc9;
mem[3231] = 8'h3a;
mem[3232] = 8'hd0;
mem[3233] = 8'hfe;
mem[3234] = 8'h28;
mem[3235] = 8'h08;
mem[3236] = 8'hca;
mem[3237] = 8'h28;
mem[3238] = 8'h8a;
mem[3239] = 8'h08;
mem[3240] = 8'hc9;
mem[3241] = 8'hff;
mem[3242] = 8'hd0;
mem[3243] = 8'hfe;
mem[3244] = 8'h68;
mem[3245] = 8'h48;
mem[3246] = 8'h09;
mem[3247] = 8'h08;
mem[3248] = 8'hc9;
mem[3249] = 8'hb8;
mem[3250] = 8'hd0;
mem[3251] = 8'hfe;
mem[3252] = 8'h28;
mem[3253] = 8'ha0;
mem[3254] = 8'hff;
mem[3255] = 8'ha9;
mem[3256] = 8'hff;
mem[3257] = 8'h48;
mem[3258] = 8'h28;
mem[3259] = 8'h98;
mem[3260] = 8'h08;
mem[3261] = 8'hc9;
mem[3262] = 8'hff;
mem[3263] = 8'hd0;
mem[3264] = 8'hfe;
mem[3265] = 8'h68;
mem[3266] = 8'h48;
mem[3267] = 8'h09;
mem[3268] = 8'h08;
mem[3269] = 8'hc9;
mem[3270] = 8'hfd;
mem[3271] = 8'hd0;
mem[3272] = 8'hfe;
mem[3273] = 8'h28;
mem[3274] = 8'h08;
mem[3275] = 8'hc8;
mem[3276] = 8'h28;
mem[3277] = 8'h98;
mem[3278] = 8'h08;
mem[3279] = 8'hc9;
mem[3280] = 8'h00;
mem[3281] = 8'hd0;
mem[3282] = 8'hfe;
mem[3283] = 8'h68;
mem[3284] = 8'h48;
mem[3285] = 8'h09;
mem[3286] = 8'h08;
mem[3287] = 8'hc9;
mem[3288] = 8'h7f;
mem[3289] = 8'hd0;
mem[3290] = 8'hfe;
mem[3291] = 8'h28;
mem[3292] = 8'h08;
mem[3293] = 8'hc8;
mem[3294] = 8'h28;
mem[3295] = 8'h98;
mem[3296] = 8'h08;
mem[3297] = 8'hc9;
mem[3298] = 8'h01;
mem[3299] = 8'hd0;
mem[3300] = 8'hfe;
mem[3301] = 8'h68;
mem[3302] = 8'h48;
mem[3303] = 8'h09;
mem[3304] = 8'h08;
mem[3305] = 8'hc9;
mem[3306] = 8'h7d;
mem[3307] = 8'hd0;
mem[3308] = 8'hfe;
mem[3309] = 8'h28;
mem[3310] = 8'ha9;
mem[3311] = 8'h00;
mem[3312] = 8'h48;
mem[3313] = 8'h28;
mem[3314] = 8'h98;
mem[3315] = 8'h08;
mem[3316] = 8'hc9;
mem[3317] = 8'h01;
mem[3318] = 8'hd0;
mem[3319] = 8'hfe;
mem[3320] = 8'h68;
mem[3321] = 8'h48;
mem[3322] = 8'h09;
mem[3323] = 8'h08;
mem[3324] = 8'hc9;
mem[3325] = 8'h38;
mem[3326] = 8'hd0;
mem[3327] = 8'hfe;
mem[3328] = 8'h28;
mem[3329] = 8'h08;
mem[3330] = 8'h88;
mem[3331] = 8'h28;
mem[3332] = 8'h98;
mem[3333] = 8'h08;
mem[3334] = 8'hc9;
mem[3335] = 8'h00;
mem[3336] = 8'hd0;
mem[3337] = 8'hfe;
mem[3338] = 8'h68;
mem[3339] = 8'h48;
mem[3340] = 8'h09;
mem[3341] = 8'h08;
mem[3342] = 8'hc9;
mem[3343] = 8'h3a;
mem[3344] = 8'hd0;
mem[3345] = 8'hfe;
mem[3346] = 8'h28;
mem[3347] = 8'h08;
mem[3348] = 8'h88;
mem[3349] = 8'h28;
mem[3350] = 8'h98;
mem[3351] = 8'h08;
mem[3352] = 8'hc9;
mem[3353] = 8'hff;
mem[3354] = 8'hd0;
mem[3355] = 8'hfe;
mem[3356] = 8'h68;
mem[3357] = 8'h48;
mem[3358] = 8'h09;
mem[3359] = 8'h08;
mem[3360] = 8'hc9;
mem[3361] = 8'hb8;
mem[3362] = 8'hd0;
mem[3363] = 8'hfe;
mem[3364] = 8'h28;
mem[3365] = 8'ha9;
mem[3366] = 8'hff;
mem[3367] = 8'h48;
mem[3368] = 8'ha2;
mem[3369] = 8'hff;
mem[3370] = 8'h8a;
mem[3371] = 8'h28;
mem[3372] = 8'ha8;
mem[3373] = 8'h08;
mem[3374] = 8'hc0;
mem[3375] = 8'hff;
mem[3376] = 8'hd0;
mem[3377] = 8'hfe;
mem[3378] = 8'h68;
mem[3379] = 8'h48;
mem[3380] = 8'h09;
mem[3381] = 8'h08;
mem[3382] = 8'hc9;
mem[3383] = 8'hfd;
mem[3384] = 8'hd0;
mem[3385] = 8'hfe;
mem[3386] = 8'h28;
mem[3387] = 8'h08;
mem[3388] = 8'he8;
mem[3389] = 8'h8a;
mem[3390] = 8'h28;
mem[3391] = 8'ha8;
mem[3392] = 8'h08;
mem[3393] = 8'hc0;
mem[3394] = 8'h00;
mem[3395] = 8'hd0;
mem[3396] = 8'hfe;
mem[3397] = 8'h68;
mem[3398] = 8'h48;
mem[3399] = 8'h09;
mem[3400] = 8'h08;
mem[3401] = 8'hc9;
mem[3402] = 8'h7f;
mem[3403] = 8'hd0;
mem[3404] = 8'hfe;
mem[3405] = 8'h28;
mem[3406] = 8'h08;
mem[3407] = 8'he8;
mem[3408] = 8'h8a;
mem[3409] = 8'h28;
mem[3410] = 8'ha8;
mem[3411] = 8'h08;
mem[3412] = 8'hc0;
mem[3413] = 8'h01;
mem[3414] = 8'hd0;
mem[3415] = 8'hfe;
mem[3416] = 8'h68;
mem[3417] = 8'h48;
mem[3418] = 8'h09;
mem[3419] = 8'h08;
mem[3420] = 8'hc9;
mem[3421] = 8'h7d;
mem[3422] = 8'hd0;
mem[3423] = 8'hfe;
mem[3424] = 8'h28;
mem[3425] = 8'ha9;
mem[3426] = 8'h00;
mem[3427] = 8'h48;
mem[3428] = 8'ha9;
mem[3429] = 8'h00;
mem[3430] = 8'h8a;
mem[3431] = 8'h28;
mem[3432] = 8'ha8;
mem[3433] = 8'h08;
mem[3434] = 8'hc0;
mem[3435] = 8'h01;
mem[3436] = 8'hd0;
mem[3437] = 8'hfe;
mem[3438] = 8'h68;
mem[3439] = 8'h48;
mem[3440] = 8'h09;
mem[3441] = 8'h08;
mem[3442] = 8'hc9;
mem[3443] = 8'h38;
mem[3444] = 8'hd0;
mem[3445] = 8'hfe;
mem[3446] = 8'h28;
mem[3447] = 8'h08;
mem[3448] = 8'hca;
mem[3449] = 8'h8a;
mem[3450] = 8'h28;
mem[3451] = 8'ha8;
mem[3452] = 8'h08;
mem[3453] = 8'hc0;
mem[3454] = 8'h00;
mem[3455] = 8'hd0;
mem[3456] = 8'hfe;
mem[3457] = 8'h68;
mem[3458] = 8'h48;
mem[3459] = 8'h09;
mem[3460] = 8'h08;
mem[3461] = 8'hc9;
mem[3462] = 8'h3a;
mem[3463] = 8'hd0;
mem[3464] = 8'hfe;
mem[3465] = 8'h28;
mem[3466] = 8'h08;
mem[3467] = 8'hca;
mem[3468] = 8'h8a;
mem[3469] = 8'h28;
mem[3470] = 8'ha8;
mem[3471] = 8'h08;
mem[3472] = 8'hc0;
mem[3473] = 8'hff;
mem[3474] = 8'hd0;
mem[3475] = 8'hfe;
mem[3476] = 8'h68;
mem[3477] = 8'h48;
mem[3478] = 8'h09;
mem[3479] = 8'h08;
mem[3480] = 8'hc9;
mem[3481] = 8'hb8;
mem[3482] = 8'hd0;
mem[3483] = 8'hfe;
mem[3484] = 8'h28;
mem[3485] = 8'ha9;
mem[3486] = 8'hff;
mem[3487] = 8'h48;
mem[3488] = 8'ha0;
mem[3489] = 8'hff;
mem[3490] = 8'h98;
mem[3491] = 8'h28;
mem[3492] = 8'haa;
mem[3493] = 8'h08;
mem[3494] = 8'he0;
mem[3495] = 8'hff;
mem[3496] = 8'hd0;
mem[3497] = 8'hfe;
mem[3498] = 8'h68;
mem[3499] = 8'h48;
mem[3500] = 8'h09;
mem[3501] = 8'h08;
mem[3502] = 8'hc9;
mem[3503] = 8'hfd;
mem[3504] = 8'hd0;
mem[3505] = 8'hfe;
mem[3506] = 8'h28;
mem[3507] = 8'h08;
mem[3508] = 8'hc8;
mem[3509] = 8'h98;
mem[3510] = 8'h28;
mem[3511] = 8'haa;
mem[3512] = 8'h08;
mem[3513] = 8'he0;
mem[3514] = 8'h00;
mem[3515] = 8'hd0;
mem[3516] = 8'hfe;
mem[3517] = 8'h68;
mem[3518] = 8'h48;
mem[3519] = 8'h09;
mem[3520] = 8'h08;
mem[3521] = 8'hc9;
mem[3522] = 8'h7f;
mem[3523] = 8'hd0;
mem[3524] = 8'hfe;
mem[3525] = 8'h28;
mem[3526] = 8'h08;
mem[3527] = 8'hc8;
mem[3528] = 8'h98;
mem[3529] = 8'h28;
mem[3530] = 8'haa;
mem[3531] = 8'h08;
mem[3532] = 8'he0;
mem[3533] = 8'h01;
mem[3534] = 8'hd0;
mem[3535] = 8'hfe;
mem[3536] = 8'h68;
mem[3537] = 8'h48;
mem[3538] = 8'h09;
mem[3539] = 8'h08;
mem[3540] = 8'hc9;
mem[3541] = 8'h7d;
mem[3542] = 8'hd0;
mem[3543] = 8'hfe;
mem[3544] = 8'h28;
mem[3545] = 8'ha9;
mem[3546] = 8'h00;
mem[3547] = 8'h48;
mem[3548] = 8'ha9;
mem[3549] = 8'h00;
mem[3550] = 8'h98;
mem[3551] = 8'h28;
mem[3552] = 8'haa;
mem[3553] = 8'h08;
mem[3554] = 8'he0;
mem[3555] = 8'h01;
mem[3556] = 8'hd0;
mem[3557] = 8'hfe;
mem[3558] = 8'h68;
mem[3559] = 8'h48;
mem[3560] = 8'h09;
mem[3561] = 8'h08;
mem[3562] = 8'hc9;
mem[3563] = 8'h38;
mem[3564] = 8'hd0;
mem[3565] = 8'hfe;
mem[3566] = 8'h28;
mem[3567] = 8'h08;
mem[3568] = 8'h88;
mem[3569] = 8'h98;
mem[3570] = 8'h28;
mem[3571] = 8'haa;
mem[3572] = 8'h08;
mem[3573] = 8'he0;
mem[3574] = 8'h00;
mem[3575] = 8'hd0;
mem[3576] = 8'hfe;
mem[3577] = 8'h68;
mem[3578] = 8'h48;
mem[3579] = 8'h09;
mem[3580] = 8'h08;
mem[3581] = 8'hc9;
mem[3582] = 8'h3a;
mem[3583] = 8'hd0;
mem[3584] = 8'hfe;
mem[3585] = 8'h28;
mem[3586] = 8'h08;
mem[3587] = 8'h88;
mem[3588] = 8'h98;
mem[3589] = 8'h28;
mem[3590] = 8'haa;
mem[3591] = 8'h08;
mem[3592] = 8'he0;
mem[3593] = 8'hff;
mem[3594] = 8'hd0;
mem[3595] = 8'hfe;
mem[3596] = 8'h68;
mem[3597] = 8'h48;
mem[3598] = 8'h09;
mem[3599] = 8'h08;
mem[3600] = 8'hc9;
mem[3601] = 8'hb8;
mem[3602] = 8'hd0;
mem[3603] = 8'hfe;
mem[3604] = 8'h28;
mem[3605] = 8'had;
mem[3606] = 8'h00;
mem[3607] = 8'h02;
mem[3608] = 8'hc9;
mem[3609] = 8'h0d;
mem[3610] = 8'hd0;
mem[3611] = 8'hfe;
mem[3612] = 8'ha9;
mem[3613] = 8'h0e;
mem[3614] = 8'h8d;
mem[3615] = 8'h00;
mem[3616] = 8'h02;
mem[3617] = 8'ha2;
mem[3618] = 8'h01;
mem[3619] = 8'ha9;
mem[3620] = 8'hff;
mem[3621] = 8'h48;
mem[3622] = 8'h28;
mem[3623] = 8'h9a;
mem[3624] = 8'h08;
mem[3625] = 8'had;
mem[3626] = 8'h01;
mem[3627] = 8'h01;
mem[3628] = 8'h09;
mem[3629] = 8'h08;
mem[3630] = 8'hc9;
mem[3631] = 8'hff;
mem[3632] = 8'hd0;
mem[3633] = 8'hfe;
mem[3634] = 8'ha9;
mem[3635] = 8'h00;
mem[3636] = 8'h48;
mem[3637] = 8'h28;
mem[3638] = 8'h9a;
mem[3639] = 8'h08;
mem[3640] = 8'had;
mem[3641] = 8'h01;
mem[3642] = 8'h01;
mem[3643] = 8'h09;
mem[3644] = 8'h08;
mem[3645] = 8'hc9;
mem[3646] = 8'h38;
mem[3647] = 8'hd0;
mem[3648] = 8'hfe;
mem[3649] = 8'hca;
mem[3650] = 8'ha9;
mem[3651] = 8'hff;
mem[3652] = 8'h48;
mem[3653] = 8'h28;
mem[3654] = 8'h9a;
mem[3655] = 8'h08;
mem[3656] = 8'had;
mem[3657] = 8'h00;
mem[3658] = 8'h01;
mem[3659] = 8'h09;
mem[3660] = 8'h08;
mem[3661] = 8'hc9;
mem[3662] = 8'hff;
mem[3663] = 8'hd0;
mem[3664] = 8'hfe;
mem[3665] = 8'ha9;
mem[3666] = 8'h00;
mem[3667] = 8'h48;
mem[3668] = 8'h28;
mem[3669] = 8'h9a;
mem[3670] = 8'h08;
mem[3671] = 8'had;
mem[3672] = 8'h00;
mem[3673] = 8'h01;
mem[3674] = 8'h09;
mem[3675] = 8'h08;
mem[3676] = 8'hc9;
mem[3677] = 8'h38;
mem[3678] = 8'hd0;
mem[3679] = 8'hfe;
mem[3680] = 8'hca;
mem[3681] = 8'ha9;
mem[3682] = 8'hff;
mem[3683] = 8'h48;
mem[3684] = 8'h28;
mem[3685] = 8'h9a;
mem[3686] = 8'h08;
mem[3687] = 8'had;
mem[3688] = 8'hff;
mem[3689] = 8'h01;
mem[3690] = 8'h09;
mem[3691] = 8'h08;
mem[3692] = 8'hc9;
mem[3693] = 8'hff;
mem[3694] = 8'hd0;
mem[3695] = 8'hfe;
mem[3696] = 8'ha9;
mem[3697] = 8'h00;
mem[3698] = 8'h48;
mem[3699] = 8'h28;
mem[3700] = 8'h9a;
mem[3701] = 8'h08;
mem[3702] = 8'had;
mem[3703] = 8'hff;
mem[3704] = 8'h01;
mem[3705] = 8'h09;
mem[3706] = 8'h08;
mem[3707] = 8'hc9;
mem[3708] = 8'h38;
mem[3709] = 8'ha2;
mem[3710] = 8'h01;
mem[3711] = 8'h9a;
mem[3712] = 8'ha9;
mem[3713] = 8'hff;
mem[3714] = 8'h48;
mem[3715] = 8'h28;
mem[3716] = 8'hba;
mem[3717] = 8'h08;
mem[3718] = 8'he0;
mem[3719] = 8'h01;
mem[3720] = 8'hd0;
mem[3721] = 8'hfe;
mem[3722] = 8'had;
mem[3723] = 8'h01;
mem[3724] = 8'h01;
mem[3725] = 8'h09;
mem[3726] = 8'h08;
mem[3727] = 8'hc9;
mem[3728] = 8'h7d;
mem[3729] = 8'hd0;
mem[3730] = 8'hfe;
mem[3731] = 8'ha9;
mem[3732] = 8'hff;
mem[3733] = 8'h48;
mem[3734] = 8'h28;
mem[3735] = 8'hba;
mem[3736] = 8'h08;
mem[3737] = 8'he0;
mem[3738] = 8'h00;
mem[3739] = 8'hd0;
mem[3740] = 8'hfe;
mem[3741] = 8'had;
mem[3742] = 8'h00;
mem[3743] = 8'h01;
mem[3744] = 8'h09;
mem[3745] = 8'h08;
mem[3746] = 8'hc9;
mem[3747] = 8'h7f;
mem[3748] = 8'hd0;
mem[3749] = 8'hfe;
mem[3750] = 8'ha9;
mem[3751] = 8'hff;
mem[3752] = 8'h48;
mem[3753] = 8'h28;
mem[3754] = 8'hba;
mem[3755] = 8'h08;
mem[3756] = 8'he0;
mem[3757] = 8'hff;
mem[3758] = 8'hd0;
mem[3759] = 8'hfe;
mem[3760] = 8'had;
mem[3761] = 8'hff;
mem[3762] = 8'h01;
mem[3763] = 8'h09;
mem[3764] = 8'h08;
mem[3765] = 8'hc9;
mem[3766] = 8'hfd;
mem[3767] = 8'hd0;
mem[3768] = 8'hfe;
mem[3769] = 8'ha2;
mem[3770] = 8'h01;
mem[3771] = 8'h9a;
mem[3772] = 8'ha9;
mem[3773] = 8'h00;
mem[3774] = 8'h48;
mem[3775] = 8'h28;
mem[3776] = 8'hba;
mem[3777] = 8'h08;
mem[3778] = 8'he0;
mem[3779] = 8'h01;
mem[3780] = 8'hd0;
mem[3781] = 8'hfe;
mem[3782] = 8'had;
mem[3783] = 8'h01;
mem[3784] = 8'h01;
mem[3785] = 8'h09;
mem[3786] = 8'h08;
mem[3787] = 8'hc9;
mem[3788] = 8'h38;
mem[3789] = 8'hd0;
mem[3790] = 8'hfe;
mem[3791] = 8'ha9;
mem[3792] = 8'h00;
mem[3793] = 8'h48;
mem[3794] = 8'h28;
mem[3795] = 8'hba;
mem[3796] = 8'h08;
mem[3797] = 8'he0;
mem[3798] = 8'h00;
mem[3799] = 8'hd0;
mem[3800] = 8'hfe;
mem[3801] = 8'had;
mem[3802] = 8'h00;
mem[3803] = 8'h01;
mem[3804] = 8'h09;
mem[3805] = 8'h08;
mem[3806] = 8'hc9;
mem[3807] = 8'h3a;
mem[3808] = 8'hd0;
mem[3809] = 8'hfe;
mem[3810] = 8'ha9;
mem[3811] = 8'h00;
mem[3812] = 8'h48;
mem[3813] = 8'h28;
mem[3814] = 8'hba;
mem[3815] = 8'h08;
mem[3816] = 8'he0;
mem[3817] = 8'hff;
mem[3818] = 8'hd0;
mem[3819] = 8'hfe;
mem[3820] = 8'had;
mem[3821] = 8'hff;
mem[3822] = 8'h01;
mem[3823] = 8'h09;
mem[3824] = 8'h08;
mem[3825] = 8'hc9;
mem[3826] = 8'hb8;
mem[3827] = 8'hd0;
mem[3828] = 8'hfe;
mem[3829] = 8'h68;
mem[3830] = 8'had;
mem[3831] = 8'h00;
mem[3832] = 8'h02;
mem[3833] = 8'hc9;
mem[3834] = 8'h0e;
mem[3835] = 8'hd0;
mem[3836] = 8'hfe;
mem[3837] = 8'ha9;
mem[3838] = 8'h0f;
mem[3839] = 8'h8d;
mem[3840] = 8'h00;
mem[3841] = 8'h02;
mem[3842] = 8'ha0;
mem[3843] = 8'h03;
mem[3844] = 8'ha9;
mem[3845] = 8'h00;
mem[3846] = 8'h48;
mem[3847] = 8'h28;
mem[3848] = 8'hb6;
mem[3849] = 8'h13;
mem[3850] = 8'h08;
mem[3851] = 8'h8a;
mem[3852] = 8'h49;
mem[3853] = 8'hc3;
mem[3854] = 8'h28;
mem[3855] = 8'h99;
mem[3856] = 8'h03;
mem[3857] = 8'h02;
mem[3858] = 8'h08;
mem[3859] = 8'h49;
mem[3860] = 8'hc3;
mem[3861] = 8'hd9;
mem[3862] = 8'h17;
mem[3863] = 8'h02;
mem[3864] = 8'hd0;
mem[3865] = 8'hfe;
mem[3866] = 8'h68;
mem[3867] = 8'h09;
mem[3868] = 8'h08;
mem[3869] = 8'h49;
mem[3870] = 8'h38;
mem[3871] = 8'hd9;
mem[3872] = 8'h1c;
mem[3873] = 8'h02;
mem[3874] = 8'hd0;
mem[3875] = 8'hfe;
mem[3876] = 8'h88;
mem[3877] = 8'h10;
mem[3878] = 8'hdd;
mem[3879] = 8'ha0;
mem[3880] = 8'h03;
mem[3881] = 8'ha9;
mem[3882] = 8'hff;
mem[3883] = 8'h48;
mem[3884] = 8'h28;
mem[3885] = 8'hb6;
mem[3886] = 8'h13;
mem[3887] = 8'h08;
mem[3888] = 8'h8a;
mem[3889] = 8'h49;
mem[3890] = 8'hc3;
mem[3891] = 8'h28;
mem[3892] = 8'h99;
mem[3893] = 8'h03;
mem[3894] = 8'h02;
mem[3895] = 8'h08;
mem[3896] = 8'h49;
mem[3897] = 8'hc3;
mem[3898] = 8'hd9;
mem[3899] = 8'h17;
mem[3900] = 8'h02;
mem[3901] = 8'hd0;
mem[3902] = 8'hfe;
mem[3903] = 8'h68;
mem[3904] = 8'h09;
mem[3905] = 8'h08;
mem[3906] = 8'h49;
mem[3907] = 8'h7d;
mem[3908] = 8'hd9;
mem[3909] = 8'h1c;
mem[3910] = 8'h02;
mem[3911] = 8'hd0;
mem[3912] = 8'hfe;
mem[3913] = 8'h88;
mem[3914] = 8'h10;
mem[3915] = 8'hdd;
mem[3916] = 8'ha0;
mem[3917] = 8'h03;
mem[3918] = 8'ha9;
mem[3919] = 8'h00;
mem[3920] = 8'h48;
mem[3921] = 8'h28;
mem[3922] = 8'hbe;
mem[3923] = 8'h17;
mem[3924] = 8'h02;
mem[3925] = 8'h08;
mem[3926] = 8'h8a;
mem[3927] = 8'h49;
mem[3928] = 8'hc3;
mem[3929] = 8'haa;
mem[3930] = 8'h28;
mem[3931] = 8'h96;
mem[3932] = 8'h0c;
mem[3933] = 8'h08;
mem[3934] = 8'h49;
mem[3935] = 8'hc3;
mem[3936] = 8'hd9;
mem[3937] = 8'h13;
mem[3938] = 8'h00;
mem[3939] = 8'hd0;
mem[3940] = 8'hfe;
mem[3941] = 8'h68;
mem[3942] = 8'h09;
mem[3943] = 8'h08;
mem[3944] = 8'h49;
mem[3945] = 8'h38;
mem[3946] = 8'hd9;
mem[3947] = 8'h1c;
mem[3948] = 8'h02;
mem[3949] = 8'hd0;
mem[3950] = 8'hfe;
mem[3951] = 8'h88;
mem[3952] = 8'h10;
mem[3953] = 8'hdc;
mem[3954] = 8'ha0;
mem[3955] = 8'h03;
mem[3956] = 8'ha9;
mem[3957] = 8'hff;
mem[3958] = 8'h48;
mem[3959] = 8'h28;
mem[3960] = 8'hbe;
mem[3961] = 8'h17;
mem[3962] = 8'h02;
mem[3963] = 8'h08;
mem[3964] = 8'h8a;
mem[3965] = 8'h49;
mem[3966] = 8'hc3;
mem[3967] = 8'haa;
mem[3968] = 8'h28;
mem[3969] = 8'h96;
mem[3970] = 8'h0c;
mem[3971] = 8'h08;
mem[3972] = 8'h49;
mem[3973] = 8'hc3;
mem[3974] = 8'hd9;
mem[3975] = 8'h13;
mem[3976] = 8'h00;
mem[3977] = 8'hd0;
mem[3978] = 8'hfe;
mem[3979] = 8'h68;
mem[3980] = 8'h09;
mem[3981] = 8'h08;
mem[3982] = 8'h49;
mem[3983] = 8'h7d;
mem[3984] = 8'hd9;
mem[3985] = 8'h1c;
mem[3986] = 8'h02;
mem[3987] = 8'hd0;
mem[3988] = 8'hfe;
mem[3989] = 8'h88;
mem[3990] = 8'h10;
mem[3991] = 8'hdc;
mem[3992] = 8'ha0;
mem[3993] = 8'h03;
mem[3994] = 8'ha2;
mem[3995] = 8'h00;
mem[3996] = 8'hb9;
mem[3997] = 8'h0c;
mem[3998] = 8'h00;
mem[3999] = 8'h49;
mem[4000] = 8'hc3;
mem[4001] = 8'hd9;
mem[4002] = 8'h13;
mem[4003] = 8'h00;
mem[4004] = 8'hd0;
mem[4005] = 8'hfe;
mem[4006] = 8'h96;
mem[4007] = 8'h0c;
mem[4008] = 8'hb9;
mem[4009] = 8'h03;
mem[4010] = 8'h02;
mem[4011] = 8'h49;
mem[4012] = 8'hc3;
mem[4013] = 8'hd9;
mem[4014] = 8'h17;
mem[4015] = 8'h02;
mem[4016] = 8'hd0;
mem[4017] = 8'hfe;
mem[4018] = 8'h8a;
mem[4019] = 8'h99;
mem[4020] = 8'h03;
mem[4021] = 8'h02;
mem[4022] = 8'h88;
mem[4023] = 8'h10;
mem[4024] = 8'he3;
mem[4025] = 8'had;
mem[4026] = 8'h00;
mem[4027] = 8'h02;
mem[4028] = 8'hc9;
mem[4029] = 8'h0f;
mem[4030] = 8'hd0;
mem[4031] = 8'hfe;
mem[4032] = 8'ha9;
mem[4033] = 8'h10;
mem[4034] = 8'h8d;
mem[4035] = 8'h00;
mem[4036] = 8'h02;
mem[4037] = 8'ha0;
mem[4038] = 8'hfd;
mem[4039] = 8'hb6;
mem[4040] = 8'h19;
mem[4041] = 8'h8a;
mem[4042] = 8'h99;
mem[4043] = 8'h09;
mem[4044] = 8'h01;
mem[4045] = 8'h88;
mem[4046] = 8'hc0;
mem[4047] = 8'hfa;
mem[4048] = 8'hb0;
mem[4049] = 8'hf5;
mem[4050] = 8'ha0;
mem[4051] = 8'hfd;
mem[4052] = 8'hbe;
mem[4053] = 8'h1d;
mem[4054] = 8'h01;
mem[4055] = 8'h96;
mem[4056] = 8'h12;
mem[4057] = 8'h88;
mem[4058] = 8'hc0;
mem[4059] = 8'hfa;
mem[4060] = 8'hb0;
mem[4061] = 8'hf6;
mem[4062] = 8'ha0;
mem[4063] = 8'h03;
mem[4064] = 8'ha2;
mem[4065] = 8'h00;
mem[4066] = 8'hb9;
mem[4067] = 8'h0c;
mem[4068] = 8'h00;
mem[4069] = 8'hd9;
mem[4070] = 8'h13;
mem[4071] = 8'h00;
mem[4072] = 8'hd0;
mem[4073] = 8'hfe;
mem[4074] = 8'h96;
mem[4075] = 8'h0c;
mem[4076] = 8'hb9;
mem[4077] = 8'h03;
mem[4078] = 8'h02;
mem[4079] = 8'hd9;
mem[4080] = 8'h17;
mem[4081] = 8'h02;
mem[4082] = 8'hd0;
mem[4083] = 8'hfe;
mem[4084] = 8'h8a;
mem[4085] = 8'h99;
mem[4086] = 8'h03;
mem[4087] = 8'h02;
mem[4088] = 8'h88;
mem[4089] = 8'h10;
mem[4090] = 8'he7;
mem[4091] = 8'had;
mem[4092] = 8'h00;
mem[4093] = 8'h02;
mem[4094] = 8'hc9;
mem[4095] = 8'h10;
mem[4096] = 8'hd0;
mem[4097] = 8'hfe;
mem[4098] = 8'ha9;
mem[4099] = 8'h11;
mem[4100] = 8'h8d;
mem[4101] = 8'h00;
mem[4102] = 8'h02;
mem[4103] = 8'ha2;
mem[4104] = 8'h03;
mem[4105] = 8'ha9;
mem[4106] = 8'h00;
mem[4107] = 8'h48;
mem[4108] = 8'h28;
mem[4109] = 8'hb4;
mem[4110] = 8'h13;
mem[4111] = 8'h08;
mem[4112] = 8'h98;
mem[4113] = 8'h49;
mem[4114] = 8'hc3;
mem[4115] = 8'h28;
mem[4116] = 8'h9d;
mem[4117] = 8'h03;
mem[4118] = 8'h02;
mem[4119] = 8'h08;
mem[4120] = 8'h49;
mem[4121] = 8'hc3;
mem[4122] = 8'hdd;
mem[4123] = 8'h17;
mem[4124] = 8'h02;
mem[4125] = 8'hd0;
mem[4126] = 8'hfe;
mem[4127] = 8'h68;
mem[4128] = 8'h09;
mem[4129] = 8'h08;
mem[4130] = 8'h49;
mem[4131] = 8'h38;
mem[4132] = 8'hdd;
mem[4133] = 8'h1c;
mem[4134] = 8'h02;
mem[4135] = 8'hd0;
mem[4136] = 8'hfe;
mem[4137] = 8'hca;
mem[4138] = 8'h10;
mem[4139] = 8'hdd;
mem[4140] = 8'ha2;
mem[4141] = 8'h03;
mem[4142] = 8'ha9;
mem[4143] = 8'hff;
mem[4144] = 8'h48;
mem[4145] = 8'h28;
mem[4146] = 8'hb4;
mem[4147] = 8'h13;
mem[4148] = 8'h08;
mem[4149] = 8'h98;
mem[4150] = 8'h49;
mem[4151] = 8'hc3;
mem[4152] = 8'h28;
mem[4153] = 8'h9d;
mem[4154] = 8'h03;
mem[4155] = 8'h02;
mem[4156] = 8'h08;
mem[4157] = 8'h49;
mem[4158] = 8'hc3;
mem[4159] = 8'hdd;
mem[4160] = 8'h17;
mem[4161] = 8'h02;
mem[4162] = 8'hd0;
mem[4163] = 8'hfe;
mem[4164] = 8'h68;
mem[4165] = 8'h09;
mem[4166] = 8'h08;
mem[4167] = 8'h49;
mem[4168] = 8'h7d;
mem[4169] = 8'hdd;
mem[4170] = 8'h1c;
mem[4171] = 8'h02;
mem[4172] = 8'hd0;
mem[4173] = 8'hfe;
mem[4174] = 8'hca;
mem[4175] = 8'h10;
mem[4176] = 8'hdd;
mem[4177] = 8'ha2;
mem[4178] = 8'h03;
mem[4179] = 8'ha9;
mem[4180] = 8'h00;
mem[4181] = 8'h48;
mem[4182] = 8'h28;
mem[4183] = 8'hbc;
mem[4184] = 8'h17;
mem[4185] = 8'h02;
mem[4186] = 8'h08;
mem[4187] = 8'h98;
mem[4188] = 8'h49;
mem[4189] = 8'hc3;
mem[4190] = 8'ha8;
mem[4191] = 8'h28;
mem[4192] = 8'h94;
mem[4193] = 8'h0c;
mem[4194] = 8'h08;
mem[4195] = 8'h49;
mem[4196] = 8'hc3;
mem[4197] = 8'hd5;
mem[4198] = 8'h13;
mem[4199] = 8'hd0;
mem[4200] = 8'hfe;
mem[4201] = 8'h68;
mem[4202] = 8'h09;
mem[4203] = 8'h08;
mem[4204] = 8'h49;
mem[4205] = 8'h38;
mem[4206] = 8'hdd;
mem[4207] = 8'h1c;
mem[4208] = 8'h02;
mem[4209] = 8'hd0;
mem[4210] = 8'hfe;
mem[4211] = 8'hca;
mem[4212] = 8'h10;
mem[4213] = 8'hdd;
mem[4214] = 8'ha2;
mem[4215] = 8'h03;
mem[4216] = 8'ha9;
mem[4217] = 8'hff;
mem[4218] = 8'h48;
mem[4219] = 8'h28;
mem[4220] = 8'hbc;
mem[4221] = 8'h17;
mem[4222] = 8'h02;
mem[4223] = 8'h08;
mem[4224] = 8'h98;
mem[4225] = 8'h49;
mem[4226] = 8'hc3;
mem[4227] = 8'ha8;
mem[4228] = 8'h28;
mem[4229] = 8'h94;
mem[4230] = 8'h0c;
mem[4231] = 8'h08;
mem[4232] = 8'h49;
mem[4233] = 8'hc3;
mem[4234] = 8'hd5;
mem[4235] = 8'h13;
mem[4236] = 8'hd0;
mem[4237] = 8'hfe;
mem[4238] = 8'h68;
mem[4239] = 8'h09;
mem[4240] = 8'h08;
mem[4241] = 8'h49;
mem[4242] = 8'h7d;
mem[4243] = 8'hdd;
mem[4244] = 8'h1c;
mem[4245] = 8'h02;
mem[4246] = 8'hd0;
mem[4247] = 8'hfe;
mem[4248] = 8'hca;
mem[4249] = 8'h10;
mem[4250] = 8'hdd;
mem[4251] = 8'ha2;
mem[4252] = 8'h03;
mem[4253] = 8'ha0;
mem[4254] = 8'h00;
mem[4255] = 8'hb5;
mem[4256] = 8'h0c;
mem[4257] = 8'h49;
mem[4258] = 8'hc3;
mem[4259] = 8'hd5;
mem[4260] = 8'h13;
mem[4261] = 8'hd0;
mem[4262] = 8'hfe;
mem[4263] = 8'h94;
mem[4264] = 8'h0c;
mem[4265] = 8'hbd;
mem[4266] = 8'h03;
mem[4267] = 8'h02;
mem[4268] = 8'h49;
mem[4269] = 8'hc3;
mem[4270] = 8'hdd;
mem[4271] = 8'h17;
mem[4272] = 8'h02;
mem[4273] = 8'hd0;
mem[4274] = 8'hfe;
mem[4275] = 8'h8a;
mem[4276] = 8'h9d;
mem[4277] = 8'h03;
mem[4278] = 8'h02;
mem[4279] = 8'hca;
mem[4280] = 8'h10;
mem[4281] = 8'he5;
mem[4282] = 8'had;
mem[4283] = 8'h00;
mem[4284] = 8'h02;
mem[4285] = 8'hc9;
mem[4286] = 8'h11;
mem[4287] = 8'hd0;
mem[4288] = 8'hfe;
mem[4289] = 8'ha9;
mem[4290] = 8'h12;
mem[4291] = 8'h8d;
mem[4292] = 8'h00;
mem[4293] = 8'h02;
mem[4294] = 8'ha2;
mem[4295] = 8'hfd;
mem[4296] = 8'hb4;
mem[4297] = 8'h19;
mem[4298] = 8'h98;
mem[4299] = 8'h9d;
mem[4300] = 8'h09;
mem[4301] = 8'h01;
mem[4302] = 8'hca;
mem[4303] = 8'he0;
mem[4304] = 8'hfa;
mem[4305] = 8'hb0;
mem[4306] = 8'hf5;
mem[4307] = 8'ha2;
mem[4308] = 8'hfd;
mem[4309] = 8'hbc;
mem[4310] = 8'h1d;
mem[4311] = 8'h01;
mem[4312] = 8'h94;
mem[4313] = 8'h12;
mem[4314] = 8'hca;
mem[4315] = 8'he0;
mem[4316] = 8'hfa;
mem[4317] = 8'hb0;
mem[4318] = 8'hf6;
mem[4319] = 8'ha2;
mem[4320] = 8'h03;
mem[4321] = 8'ha0;
mem[4322] = 8'h00;
mem[4323] = 8'hb5;
mem[4324] = 8'h0c;
mem[4325] = 8'hd5;
mem[4326] = 8'h13;
mem[4327] = 8'hd0;
mem[4328] = 8'hfe;
mem[4329] = 8'h94;
mem[4330] = 8'h0c;
mem[4331] = 8'hbd;
mem[4332] = 8'h03;
mem[4333] = 8'h02;
mem[4334] = 8'hdd;
mem[4335] = 8'h17;
mem[4336] = 8'h02;
mem[4337] = 8'hd0;
mem[4338] = 8'hfe;
mem[4339] = 8'h8a;
mem[4340] = 8'h9d;
mem[4341] = 8'h03;
mem[4342] = 8'h02;
mem[4343] = 8'hca;
mem[4344] = 8'h10;
mem[4345] = 8'he9;
mem[4346] = 8'had;
mem[4347] = 8'h00;
mem[4348] = 8'h02;
mem[4349] = 8'hc9;
mem[4350] = 8'h12;
mem[4351] = 8'hd0;
mem[4352] = 8'hfe;
mem[4353] = 8'ha9;
mem[4354] = 8'h13;
mem[4355] = 8'h8d;
mem[4356] = 8'h00;
mem[4357] = 8'h02;
mem[4358] = 8'ha9;
mem[4359] = 8'h00;
mem[4360] = 8'h48;
mem[4361] = 8'h28;
mem[4362] = 8'ha6;
mem[4363] = 8'h13;
mem[4364] = 8'h08;
mem[4365] = 8'h8a;
mem[4366] = 8'h49;
mem[4367] = 8'hc3;
mem[4368] = 8'haa;
mem[4369] = 8'h28;
mem[4370] = 8'h8e;
mem[4371] = 8'h03;
mem[4372] = 8'h02;
mem[4373] = 8'h08;
mem[4374] = 8'h49;
mem[4375] = 8'hc3;
mem[4376] = 8'haa;
mem[4377] = 8'he0;
mem[4378] = 8'hc3;
mem[4379] = 8'hd0;
mem[4380] = 8'hfe;
mem[4381] = 8'h68;
mem[4382] = 8'h09;
mem[4383] = 8'h08;
mem[4384] = 8'h49;
mem[4385] = 8'h38;
mem[4386] = 8'hcd;
mem[4387] = 8'h1c;
mem[4388] = 8'h02;
mem[4389] = 8'hd0;
mem[4390] = 8'hfe;
mem[4391] = 8'ha9;
mem[4392] = 8'h00;
mem[4393] = 8'h48;
mem[4394] = 8'h28;
mem[4395] = 8'ha6;
mem[4396] = 8'h14;
mem[4397] = 8'h08;
mem[4398] = 8'h8a;
mem[4399] = 8'h49;
mem[4400] = 8'hc3;
mem[4401] = 8'haa;
mem[4402] = 8'h28;
mem[4403] = 8'h8e;
mem[4404] = 8'h04;
mem[4405] = 8'h02;
mem[4406] = 8'h08;
mem[4407] = 8'h49;
mem[4408] = 8'hc3;
mem[4409] = 8'haa;
mem[4410] = 8'he0;
mem[4411] = 8'h82;
mem[4412] = 8'hd0;
mem[4413] = 8'hfe;
mem[4414] = 8'h68;
mem[4415] = 8'h09;
mem[4416] = 8'h08;
mem[4417] = 8'h49;
mem[4418] = 8'h38;
mem[4419] = 8'hcd;
mem[4420] = 8'h1d;
mem[4421] = 8'h02;
mem[4422] = 8'hd0;
mem[4423] = 8'hfe;
mem[4424] = 8'ha9;
mem[4425] = 8'h00;
mem[4426] = 8'h48;
mem[4427] = 8'h28;
mem[4428] = 8'ha6;
mem[4429] = 8'h15;
mem[4430] = 8'h08;
mem[4431] = 8'h8a;
mem[4432] = 8'h49;
mem[4433] = 8'hc3;
mem[4434] = 8'haa;
mem[4435] = 8'h28;
mem[4436] = 8'h8e;
mem[4437] = 8'h05;
mem[4438] = 8'h02;
mem[4439] = 8'h08;
mem[4440] = 8'h49;
mem[4441] = 8'hc3;
mem[4442] = 8'haa;
mem[4443] = 8'he0;
mem[4444] = 8'h41;
mem[4445] = 8'hd0;
mem[4446] = 8'hfe;
mem[4447] = 8'h68;
mem[4448] = 8'h09;
mem[4449] = 8'h08;
mem[4450] = 8'h49;
mem[4451] = 8'h38;
mem[4452] = 8'hcd;
mem[4453] = 8'h1e;
mem[4454] = 8'h02;
mem[4455] = 8'hd0;
mem[4456] = 8'hfe;
mem[4457] = 8'ha9;
mem[4458] = 8'h00;
mem[4459] = 8'h48;
mem[4460] = 8'h28;
mem[4461] = 8'ha6;
mem[4462] = 8'h16;
mem[4463] = 8'h08;
mem[4464] = 8'h8a;
mem[4465] = 8'h49;
mem[4466] = 8'hc3;
mem[4467] = 8'haa;
mem[4468] = 8'h28;
mem[4469] = 8'h8e;
mem[4470] = 8'h06;
mem[4471] = 8'h02;
mem[4472] = 8'h08;
mem[4473] = 8'h49;
mem[4474] = 8'hc3;
mem[4475] = 8'haa;
mem[4476] = 8'he0;
mem[4477] = 8'h00;
mem[4478] = 8'hd0;
mem[4479] = 8'hfe;
mem[4480] = 8'h68;
mem[4481] = 8'h09;
mem[4482] = 8'h08;
mem[4483] = 8'h49;
mem[4484] = 8'h38;
mem[4485] = 8'hcd;
mem[4486] = 8'h1f;
mem[4487] = 8'h02;
mem[4488] = 8'hd0;
mem[4489] = 8'hfe;
mem[4490] = 8'ha9;
mem[4491] = 8'hff;
mem[4492] = 8'h48;
mem[4493] = 8'h28;
mem[4494] = 8'ha6;
mem[4495] = 8'h13;
mem[4496] = 8'h08;
mem[4497] = 8'h8a;
mem[4498] = 8'h49;
mem[4499] = 8'hc3;
mem[4500] = 8'haa;
mem[4501] = 8'h28;
mem[4502] = 8'h8e;
mem[4503] = 8'h03;
mem[4504] = 8'h02;
mem[4505] = 8'h08;
mem[4506] = 8'h49;
mem[4507] = 8'hc3;
mem[4508] = 8'haa;
mem[4509] = 8'he0;
mem[4510] = 8'hc3;
mem[4511] = 8'hd0;
mem[4512] = 8'hfe;
mem[4513] = 8'h68;
mem[4514] = 8'h09;
mem[4515] = 8'h08;
mem[4516] = 8'h49;
mem[4517] = 8'h7d;
mem[4518] = 8'hcd;
mem[4519] = 8'h1c;
mem[4520] = 8'h02;
mem[4521] = 8'hd0;
mem[4522] = 8'hfe;
mem[4523] = 8'ha9;
mem[4524] = 8'hff;
mem[4525] = 8'h48;
mem[4526] = 8'h28;
mem[4527] = 8'ha6;
mem[4528] = 8'h14;
mem[4529] = 8'h08;
mem[4530] = 8'h8a;
mem[4531] = 8'h49;
mem[4532] = 8'hc3;
mem[4533] = 8'haa;
mem[4534] = 8'h28;
mem[4535] = 8'h8e;
mem[4536] = 8'h04;
mem[4537] = 8'h02;
mem[4538] = 8'h08;
mem[4539] = 8'h49;
mem[4540] = 8'hc3;
mem[4541] = 8'haa;
mem[4542] = 8'he0;
mem[4543] = 8'h82;
mem[4544] = 8'hd0;
mem[4545] = 8'hfe;
mem[4546] = 8'h68;
mem[4547] = 8'h09;
mem[4548] = 8'h08;
mem[4549] = 8'h49;
mem[4550] = 8'h7d;
mem[4551] = 8'hcd;
mem[4552] = 8'h1d;
mem[4553] = 8'h02;
mem[4554] = 8'hd0;
mem[4555] = 8'hfe;
mem[4556] = 8'ha9;
mem[4557] = 8'hff;
mem[4558] = 8'h48;
mem[4559] = 8'h28;
mem[4560] = 8'ha6;
mem[4561] = 8'h15;
mem[4562] = 8'h08;
mem[4563] = 8'h8a;
mem[4564] = 8'h49;
mem[4565] = 8'hc3;
mem[4566] = 8'haa;
mem[4567] = 8'h28;
mem[4568] = 8'h8e;
mem[4569] = 8'h05;
mem[4570] = 8'h02;
mem[4571] = 8'h08;
mem[4572] = 8'h49;
mem[4573] = 8'hc3;
mem[4574] = 8'haa;
mem[4575] = 8'he0;
mem[4576] = 8'h41;
mem[4577] = 8'hd0;
mem[4578] = 8'hfe;
mem[4579] = 8'h68;
mem[4580] = 8'h09;
mem[4581] = 8'h08;
mem[4582] = 8'h49;
mem[4583] = 8'h7d;
mem[4584] = 8'hcd;
mem[4585] = 8'h1e;
mem[4586] = 8'h02;
mem[4587] = 8'hd0;
mem[4588] = 8'hfe;
mem[4589] = 8'ha9;
mem[4590] = 8'hff;
mem[4591] = 8'h48;
mem[4592] = 8'h28;
mem[4593] = 8'ha6;
mem[4594] = 8'h16;
mem[4595] = 8'h08;
mem[4596] = 8'h8a;
mem[4597] = 8'h49;
mem[4598] = 8'hc3;
mem[4599] = 8'haa;
mem[4600] = 8'h28;
mem[4601] = 8'h8e;
mem[4602] = 8'h06;
mem[4603] = 8'h02;
mem[4604] = 8'h08;
mem[4605] = 8'h49;
mem[4606] = 8'hc3;
mem[4607] = 8'haa;
mem[4608] = 8'he0;
mem[4609] = 8'h00;
mem[4610] = 8'hd0;
mem[4611] = 8'hfe;
mem[4612] = 8'h68;
mem[4613] = 8'h09;
mem[4614] = 8'h08;
mem[4615] = 8'h49;
mem[4616] = 8'h7d;
mem[4617] = 8'hcd;
mem[4618] = 8'h1f;
mem[4619] = 8'h02;
mem[4620] = 8'hd0;
mem[4621] = 8'hfe;
mem[4622] = 8'ha9;
mem[4623] = 8'h00;
mem[4624] = 8'h48;
mem[4625] = 8'h28;
mem[4626] = 8'hae;
mem[4627] = 8'h17;
mem[4628] = 8'h02;
mem[4629] = 8'h08;
mem[4630] = 8'h8a;
mem[4631] = 8'h49;
mem[4632] = 8'hc3;
mem[4633] = 8'haa;
mem[4634] = 8'h28;
mem[4635] = 8'h86;
mem[4636] = 8'h0c;
mem[4637] = 8'h08;
mem[4638] = 8'h49;
mem[4639] = 8'hc3;
mem[4640] = 8'hc5;
mem[4641] = 8'h13;
mem[4642] = 8'hd0;
mem[4643] = 8'hfe;
mem[4644] = 8'h68;
mem[4645] = 8'h09;
mem[4646] = 8'h08;
mem[4647] = 8'h49;
mem[4648] = 8'h38;
mem[4649] = 8'hcd;
mem[4650] = 8'h1c;
mem[4651] = 8'h02;
mem[4652] = 8'hd0;
mem[4653] = 8'hfe;
mem[4654] = 8'ha9;
mem[4655] = 8'h00;
mem[4656] = 8'h48;
mem[4657] = 8'h28;
mem[4658] = 8'hae;
mem[4659] = 8'h18;
mem[4660] = 8'h02;
mem[4661] = 8'h08;
mem[4662] = 8'h8a;
mem[4663] = 8'h49;
mem[4664] = 8'hc3;
mem[4665] = 8'haa;
mem[4666] = 8'h28;
mem[4667] = 8'h86;
mem[4668] = 8'h0d;
mem[4669] = 8'h08;
mem[4670] = 8'h49;
mem[4671] = 8'hc3;
mem[4672] = 8'hc5;
mem[4673] = 8'h14;
mem[4674] = 8'hd0;
mem[4675] = 8'hfe;
mem[4676] = 8'h68;
mem[4677] = 8'h09;
mem[4678] = 8'h08;
mem[4679] = 8'h49;
mem[4680] = 8'h38;
mem[4681] = 8'hcd;
mem[4682] = 8'h1d;
mem[4683] = 8'h02;
mem[4684] = 8'hd0;
mem[4685] = 8'hfe;
mem[4686] = 8'ha9;
mem[4687] = 8'h00;
mem[4688] = 8'h48;
mem[4689] = 8'h28;
mem[4690] = 8'hae;
mem[4691] = 8'h19;
mem[4692] = 8'h02;
mem[4693] = 8'h08;
mem[4694] = 8'h8a;
mem[4695] = 8'h49;
mem[4696] = 8'hc3;
mem[4697] = 8'haa;
mem[4698] = 8'h28;
mem[4699] = 8'h86;
mem[4700] = 8'h0e;
mem[4701] = 8'h08;
mem[4702] = 8'h49;
mem[4703] = 8'hc3;
mem[4704] = 8'hc5;
mem[4705] = 8'h15;
mem[4706] = 8'hd0;
mem[4707] = 8'hfe;
mem[4708] = 8'h68;
mem[4709] = 8'h09;
mem[4710] = 8'h08;
mem[4711] = 8'h49;
mem[4712] = 8'h38;
mem[4713] = 8'hcd;
mem[4714] = 8'h1e;
mem[4715] = 8'h02;
mem[4716] = 8'hd0;
mem[4717] = 8'hfe;
mem[4718] = 8'ha9;
mem[4719] = 8'h00;
mem[4720] = 8'h48;
mem[4721] = 8'h28;
mem[4722] = 8'hae;
mem[4723] = 8'h1a;
mem[4724] = 8'h02;
mem[4725] = 8'h08;
mem[4726] = 8'h8a;
mem[4727] = 8'h49;
mem[4728] = 8'hc3;
mem[4729] = 8'haa;
mem[4730] = 8'h28;
mem[4731] = 8'h86;
mem[4732] = 8'h0f;
mem[4733] = 8'h08;
mem[4734] = 8'h49;
mem[4735] = 8'hc3;
mem[4736] = 8'hc5;
mem[4737] = 8'h16;
mem[4738] = 8'hd0;
mem[4739] = 8'hfe;
mem[4740] = 8'h68;
mem[4741] = 8'h09;
mem[4742] = 8'h08;
mem[4743] = 8'h49;
mem[4744] = 8'h38;
mem[4745] = 8'hcd;
mem[4746] = 8'h1f;
mem[4747] = 8'h02;
mem[4748] = 8'hd0;
mem[4749] = 8'hfe;
mem[4750] = 8'ha9;
mem[4751] = 8'hff;
mem[4752] = 8'h48;
mem[4753] = 8'h28;
mem[4754] = 8'hae;
mem[4755] = 8'h17;
mem[4756] = 8'h02;
mem[4757] = 8'h08;
mem[4758] = 8'h8a;
mem[4759] = 8'h49;
mem[4760] = 8'hc3;
mem[4761] = 8'haa;
mem[4762] = 8'h28;
mem[4763] = 8'h86;
mem[4764] = 8'h0c;
mem[4765] = 8'h08;
mem[4766] = 8'h49;
mem[4767] = 8'hc3;
mem[4768] = 8'haa;
mem[4769] = 8'he4;
mem[4770] = 8'h13;
mem[4771] = 8'hd0;
mem[4772] = 8'hfe;
mem[4773] = 8'h68;
mem[4774] = 8'h09;
mem[4775] = 8'h08;
mem[4776] = 8'h49;
mem[4777] = 8'h7d;
mem[4778] = 8'hcd;
mem[4779] = 8'h1c;
mem[4780] = 8'h02;
mem[4781] = 8'hd0;
mem[4782] = 8'hfe;
mem[4783] = 8'ha9;
mem[4784] = 8'hff;
mem[4785] = 8'h48;
mem[4786] = 8'h28;
mem[4787] = 8'hae;
mem[4788] = 8'h18;
mem[4789] = 8'h02;
mem[4790] = 8'h08;
mem[4791] = 8'h8a;
mem[4792] = 8'h49;
mem[4793] = 8'hc3;
mem[4794] = 8'haa;
mem[4795] = 8'h28;
mem[4796] = 8'h86;
mem[4797] = 8'h0d;
mem[4798] = 8'h08;
mem[4799] = 8'h49;
mem[4800] = 8'hc3;
mem[4801] = 8'haa;
mem[4802] = 8'he4;
mem[4803] = 8'h14;
mem[4804] = 8'hd0;
mem[4805] = 8'hfe;
mem[4806] = 8'h68;
mem[4807] = 8'h09;
mem[4808] = 8'h08;
mem[4809] = 8'h49;
mem[4810] = 8'h7d;
mem[4811] = 8'hcd;
mem[4812] = 8'h1d;
mem[4813] = 8'h02;
mem[4814] = 8'hd0;
mem[4815] = 8'hfe;
mem[4816] = 8'ha9;
mem[4817] = 8'hff;
mem[4818] = 8'h48;
mem[4819] = 8'h28;
mem[4820] = 8'hae;
mem[4821] = 8'h19;
mem[4822] = 8'h02;
mem[4823] = 8'h08;
mem[4824] = 8'h8a;
mem[4825] = 8'h49;
mem[4826] = 8'hc3;
mem[4827] = 8'haa;
mem[4828] = 8'h28;
mem[4829] = 8'h86;
mem[4830] = 8'h0e;
mem[4831] = 8'h08;
mem[4832] = 8'h49;
mem[4833] = 8'hc3;
mem[4834] = 8'haa;
mem[4835] = 8'he4;
mem[4836] = 8'h15;
mem[4837] = 8'hd0;
mem[4838] = 8'hfe;
mem[4839] = 8'h68;
mem[4840] = 8'h09;
mem[4841] = 8'h08;
mem[4842] = 8'h49;
mem[4843] = 8'h7d;
mem[4844] = 8'hcd;
mem[4845] = 8'h1e;
mem[4846] = 8'h02;
mem[4847] = 8'hd0;
mem[4848] = 8'hfe;
mem[4849] = 8'ha9;
mem[4850] = 8'hff;
mem[4851] = 8'h48;
mem[4852] = 8'h28;
mem[4853] = 8'hae;
mem[4854] = 8'h1a;
mem[4855] = 8'h02;
mem[4856] = 8'h08;
mem[4857] = 8'h8a;
mem[4858] = 8'h49;
mem[4859] = 8'hc3;
mem[4860] = 8'haa;
mem[4861] = 8'h28;
mem[4862] = 8'h86;
mem[4863] = 8'h0f;
mem[4864] = 8'h08;
mem[4865] = 8'h49;
mem[4866] = 8'hc3;
mem[4867] = 8'haa;
mem[4868] = 8'he4;
mem[4869] = 8'h16;
mem[4870] = 8'hd0;
mem[4871] = 8'hfe;
mem[4872] = 8'h68;
mem[4873] = 8'h09;
mem[4874] = 8'h08;
mem[4875] = 8'h49;
mem[4876] = 8'h7d;
mem[4877] = 8'hcd;
mem[4878] = 8'h1f;
mem[4879] = 8'h02;
mem[4880] = 8'hd0;
mem[4881] = 8'hfe;
mem[4882] = 8'ha9;
mem[4883] = 8'h00;
mem[4884] = 8'h48;
mem[4885] = 8'h28;
mem[4886] = 8'ha2;
mem[4887] = 8'hc3;
mem[4888] = 8'h08;
mem[4889] = 8'hec;
mem[4890] = 8'h17;
mem[4891] = 8'h02;
mem[4892] = 8'hd0;
mem[4893] = 8'hfe;
mem[4894] = 8'h68;
mem[4895] = 8'h09;
mem[4896] = 8'h08;
mem[4897] = 8'h49;
mem[4898] = 8'h38;
mem[4899] = 8'hcd;
mem[4900] = 8'h1c;
mem[4901] = 8'h02;
mem[4902] = 8'hd0;
mem[4903] = 8'hfe;
mem[4904] = 8'ha9;
mem[4905] = 8'h00;
mem[4906] = 8'h48;
mem[4907] = 8'h28;
mem[4908] = 8'ha2;
mem[4909] = 8'h82;
mem[4910] = 8'h08;
mem[4911] = 8'hec;
mem[4912] = 8'h18;
mem[4913] = 8'h02;
mem[4914] = 8'hd0;
mem[4915] = 8'hfe;
mem[4916] = 8'h68;
mem[4917] = 8'h09;
mem[4918] = 8'h08;
mem[4919] = 8'h49;
mem[4920] = 8'h38;
mem[4921] = 8'hcd;
mem[4922] = 8'h1d;
mem[4923] = 8'h02;
mem[4924] = 8'hd0;
mem[4925] = 8'hfe;
mem[4926] = 8'ha9;
mem[4927] = 8'h00;
mem[4928] = 8'h48;
mem[4929] = 8'h28;
mem[4930] = 8'ha2;
mem[4931] = 8'h41;
mem[4932] = 8'h08;
mem[4933] = 8'hec;
mem[4934] = 8'h19;
mem[4935] = 8'h02;
mem[4936] = 8'hd0;
mem[4937] = 8'hfe;
mem[4938] = 8'h68;
mem[4939] = 8'h09;
mem[4940] = 8'h08;
mem[4941] = 8'h49;
mem[4942] = 8'h38;
mem[4943] = 8'hcd;
mem[4944] = 8'h1e;
mem[4945] = 8'h02;
mem[4946] = 8'hd0;
mem[4947] = 8'hfe;
mem[4948] = 8'ha9;
mem[4949] = 8'h00;
mem[4950] = 8'h48;
mem[4951] = 8'h28;
mem[4952] = 8'ha2;
mem[4953] = 8'h00;
mem[4954] = 8'h08;
mem[4955] = 8'hec;
mem[4956] = 8'h1a;
mem[4957] = 8'h02;
mem[4958] = 8'hd0;
mem[4959] = 8'hfe;
mem[4960] = 8'h68;
mem[4961] = 8'h09;
mem[4962] = 8'h08;
mem[4963] = 8'h49;
mem[4964] = 8'h38;
mem[4965] = 8'hcd;
mem[4966] = 8'h1f;
mem[4967] = 8'h02;
mem[4968] = 8'hd0;
mem[4969] = 8'hfe;
mem[4970] = 8'ha9;
mem[4971] = 8'hff;
mem[4972] = 8'h48;
mem[4973] = 8'h28;
mem[4974] = 8'ha2;
mem[4975] = 8'hc3;
mem[4976] = 8'h08;
mem[4977] = 8'hec;
mem[4978] = 8'h17;
mem[4979] = 8'h02;
mem[4980] = 8'hd0;
mem[4981] = 8'hfe;
mem[4982] = 8'h68;
mem[4983] = 8'h09;
mem[4984] = 8'h08;
mem[4985] = 8'h49;
mem[4986] = 8'h7d;
mem[4987] = 8'hcd;
mem[4988] = 8'h1c;
mem[4989] = 8'h02;
mem[4990] = 8'hd0;
mem[4991] = 8'hfe;
mem[4992] = 8'ha9;
mem[4993] = 8'hff;
mem[4994] = 8'h48;
mem[4995] = 8'h28;
mem[4996] = 8'ha2;
mem[4997] = 8'h82;
mem[4998] = 8'h08;
mem[4999] = 8'hec;
mem[5000] = 8'h18;
mem[5001] = 8'h02;
mem[5002] = 8'hd0;
mem[5003] = 8'hfe;
mem[5004] = 8'h68;
mem[5005] = 8'h09;
mem[5006] = 8'h08;
mem[5007] = 8'h49;
mem[5008] = 8'h7d;
mem[5009] = 8'hcd;
mem[5010] = 8'h1d;
mem[5011] = 8'h02;
mem[5012] = 8'hd0;
mem[5013] = 8'hfe;
mem[5014] = 8'ha9;
mem[5015] = 8'hff;
mem[5016] = 8'h48;
mem[5017] = 8'h28;
mem[5018] = 8'ha2;
mem[5019] = 8'h41;
mem[5020] = 8'h08;
mem[5021] = 8'hec;
mem[5022] = 8'h19;
mem[5023] = 8'h02;
mem[5024] = 8'hd0;
mem[5025] = 8'hfe;
mem[5026] = 8'h68;
mem[5027] = 8'h09;
mem[5028] = 8'h08;
mem[5029] = 8'h49;
mem[5030] = 8'h7d;
mem[5031] = 8'hcd;
mem[5032] = 8'h1e;
mem[5033] = 8'h02;
mem[5034] = 8'hd0;
mem[5035] = 8'hfe;
mem[5036] = 8'ha9;
mem[5037] = 8'hff;
mem[5038] = 8'h48;
mem[5039] = 8'h28;
mem[5040] = 8'ha2;
mem[5041] = 8'h00;
mem[5042] = 8'h08;
mem[5043] = 8'hec;
mem[5044] = 8'h1a;
mem[5045] = 8'h02;
mem[5046] = 8'hd0;
mem[5047] = 8'hfe;
mem[5048] = 8'h68;
mem[5049] = 8'h09;
mem[5050] = 8'h08;
mem[5051] = 8'h49;
mem[5052] = 8'h7d;
mem[5053] = 8'hcd;
mem[5054] = 8'h1f;
mem[5055] = 8'h02;
mem[5056] = 8'hd0;
mem[5057] = 8'hfe;
mem[5058] = 8'ha2;
mem[5059] = 8'h00;
mem[5060] = 8'ha5;
mem[5061] = 8'h0c;
mem[5062] = 8'h49;
mem[5063] = 8'hc3;
mem[5064] = 8'hc5;
mem[5065] = 8'h13;
mem[5066] = 8'hd0;
mem[5067] = 8'hfe;
mem[5068] = 8'h86;
mem[5069] = 8'h0c;
mem[5070] = 8'had;
mem[5071] = 8'h03;
mem[5072] = 8'h02;
mem[5073] = 8'h49;
mem[5074] = 8'hc3;
mem[5075] = 8'hcd;
mem[5076] = 8'h17;
mem[5077] = 8'h02;
mem[5078] = 8'hd0;
mem[5079] = 8'hfe;
mem[5080] = 8'h8e;
mem[5081] = 8'h03;
mem[5082] = 8'h02;
mem[5083] = 8'ha5;
mem[5084] = 8'h0d;
mem[5085] = 8'h49;
mem[5086] = 8'hc3;
mem[5087] = 8'hc5;
mem[5088] = 8'h14;
mem[5089] = 8'hd0;
mem[5090] = 8'hfe;
mem[5091] = 8'h86;
mem[5092] = 8'h0d;
mem[5093] = 8'had;
mem[5094] = 8'h04;
mem[5095] = 8'h02;
mem[5096] = 8'h49;
mem[5097] = 8'hc3;
mem[5098] = 8'hcd;
mem[5099] = 8'h18;
mem[5100] = 8'h02;
mem[5101] = 8'hd0;
mem[5102] = 8'hfe;
mem[5103] = 8'h8e;
mem[5104] = 8'h04;
mem[5105] = 8'h02;
mem[5106] = 8'ha5;
mem[5107] = 8'h0e;
mem[5108] = 8'h49;
mem[5109] = 8'hc3;
mem[5110] = 8'hc5;
mem[5111] = 8'h15;
mem[5112] = 8'hd0;
mem[5113] = 8'hfe;
mem[5114] = 8'h86;
mem[5115] = 8'h0e;
mem[5116] = 8'had;
mem[5117] = 8'h05;
mem[5118] = 8'h02;
mem[5119] = 8'h49;
mem[5120] = 8'hc3;
mem[5121] = 8'hcd;
mem[5122] = 8'h19;
mem[5123] = 8'h02;
mem[5124] = 8'hd0;
mem[5125] = 8'hfe;
mem[5126] = 8'h8e;
mem[5127] = 8'h05;
mem[5128] = 8'h02;
mem[5129] = 8'ha5;
mem[5130] = 8'h0f;
mem[5131] = 8'h49;
mem[5132] = 8'hc3;
mem[5133] = 8'hc5;
mem[5134] = 8'h16;
mem[5135] = 8'hd0;
mem[5136] = 8'hfe;
mem[5137] = 8'h86;
mem[5138] = 8'h0f;
mem[5139] = 8'had;
mem[5140] = 8'h06;
mem[5141] = 8'h02;
mem[5142] = 8'h49;
mem[5143] = 8'hc3;
mem[5144] = 8'hcd;
mem[5145] = 8'h1a;
mem[5146] = 8'h02;
mem[5147] = 8'hd0;
mem[5148] = 8'hfe;
mem[5149] = 8'h8e;
mem[5150] = 8'h06;
mem[5151] = 8'h02;
mem[5152] = 8'had;
mem[5153] = 8'h00;
mem[5154] = 8'h02;
mem[5155] = 8'hc9;
mem[5156] = 8'h13;
mem[5157] = 8'hd0;
mem[5158] = 8'hfe;
mem[5159] = 8'ha9;
mem[5160] = 8'h14;
mem[5161] = 8'h8d;
mem[5162] = 8'h00;
mem[5163] = 8'h02;
mem[5164] = 8'ha9;
mem[5165] = 8'h00;
mem[5166] = 8'h48;
mem[5167] = 8'h28;
mem[5168] = 8'ha4;
mem[5169] = 8'h13;
mem[5170] = 8'h08;
mem[5171] = 8'h98;
mem[5172] = 8'h49;
mem[5173] = 8'hc3;
mem[5174] = 8'ha8;
mem[5175] = 8'h28;
mem[5176] = 8'h8c;
mem[5177] = 8'h03;
mem[5178] = 8'h02;
mem[5179] = 8'h08;
mem[5180] = 8'h49;
mem[5181] = 8'hc3;
mem[5182] = 8'ha8;
mem[5183] = 8'hc0;
mem[5184] = 8'hc3;
mem[5185] = 8'hd0;
mem[5186] = 8'hfe;
mem[5187] = 8'h68;
mem[5188] = 8'h09;
mem[5189] = 8'h08;
mem[5190] = 8'h49;
mem[5191] = 8'h38;
mem[5192] = 8'hcd;
mem[5193] = 8'h1c;
mem[5194] = 8'h02;
mem[5195] = 8'hd0;
mem[5196] = 8'hfe;
mem[5197] = 8'ha9;
mem[5198] = 8'h00;
mem[5199] = 8'h48;
mem[5200] = 8'h28;
mem[5201] = 8'ha4;
mem[5202] = 8'h14;
mem[5203] = 8'h08;
mem[5204] = 8'h98;
mem[5205] = 8'h49;
mem[5206] = 8'hc3;
mem[5207] = 8'ha8;
mem[5208] = 8'h28;
mem[5209] = 8'h8c;
mem[5210] = 8'h04;
mem[5211] = 8'h02;
mem[5212] = 8'h08;
mem[5213] = 8'h49;
mem[5214] = 8'hc3;
mem[5215] = 8'ha8;
mem[5216] = 8'hc0;
mem[5217] = 8'h82;
mem[5218] = 8'hd0;
mem[5219] = 8'hfe;
mem[5220] = 8'h68;
mem[5221] = 8'h09;
mem[5222] = 8'h08;
mem[5223] = 8'h49;
mem[5224] = 8'h38;
mem[5225] = 8'hcd;
mem[5226] = 8'h1d;
mem[5227] = 8'h02;
mem[5228] = 8'hd0;
mem[5229] = 8'hfe;
mem[5230] = 8'ha9;
mem[5231] = 8'h00;
mem[5232] = 8'h48;
mem[5233] = 8'h28;
mem[5234] = 8'ha4;
mem[5235] = 8'h15;
mem[5236] = 8'h08;
mem[5237] = 8'h98;
mem[5238] = 8'h49;
mem[5239] = 8'hc3;
mem[5240] = 8'ha8;
mem[5241] = 8'h28;
mem[5242] = 8'h8c;
mem[5243] = 8'h05;
mem[5244] = 8'h02;
mem[5245] = 8'h08;
mem[5246] = 8'h49;
mem[5247] = 8'hc3;
mem[5248] = 8'ha8;
mem[5249] = 8'hc0;
mem[5250] = 8'h41;
mem[5251] = 8'hd0;
mem[5252] = 8'hfe;
mem[5253] = 8'h68;
mem[5254] = 8'h09;
mem[5255] = 8'h08;
mem[5256] = 8'h49;
mem[5257] = 8'h38;
mem[5258] = 8'hcd;
mem[5259] = 8'h1e;
mem[5260] = 8'h02;
mem[5261] = 8'hd0;
mem[5262] = 8'hfe;
mem[5263] = 8'ha9;
mem[5264] = 8'h00;
mem[5265] = 8'h48;
mem[5266] = 8'h28;
mem[5267] = 8'ha4;
mem[5268] = 8'h16;
mem[5269] = 8'h08;
mem[5270] = 8'h98;
mem[5271] = 8'h49;
mem[5272] = 8'hc3;
mem[5273] = 8'ha8;
mem[5274] = 8'h28;
mem[5275] = 8'h8c;
mem[5276] = 8'h06;
mem[5277] = 8'h02;
mem[5278] = 8'h08;
mem[5279] = 8'h49;
mem[5280] = 8'hc3;
mem[5281] = 8'ha8;
mem[5282] = 8'hc0;
mem[5283] = 8'h00;
mem[5284] = 8'hd0;
mem[5285] = 8'hfe;
mem[5286] = 8'h68;
mem[5287] = 8'h09;
mem[5288] = 8'h08;
mem[5289] = 8'h49;
mem[5290] = 8'h38;
mem[5291] = 8'hcd;
mem[5292] = 8'h1f;
mem[5293] = 8'h02;
mem[5294] = 8'hd0;
mem[5295] = 8'hfe;
mem[5296] = 8'ha9;
mem[5297] = 8'hff;
mem[5298] = 8'h48;
mem[5299] = 8'h28;
mem[5300] = 8'ha4;
mem[5301] = 8'h13;
mem[5302] = 8'h08;
mem[5303] = 8'h98;
mem[5304] = 8'h49;
mem[5305] = 8'hc3;
mem[5306] = 8'ha8;
mem[5307] = 8'h28;
mem[5308] = 8'h8c;
mem[5309] = 8'h03;
mem[5310] = 8'h02;
mem[5311] = 8'h08;
mem[5312] = 8'h49;
mem[5313] = 8'hc3;
mem[5314] = 8'ha8;
mem[5315] = 8'hc0;
mem[5316] = 8'hc3;
mem[5317] = 8'hd0;
mem[5318] = 8'hfe;
mem[5319] = 8'h68;
mem[5320] = 8'h09;
mem[5321] = 8'h08;
mem[5322] = 8'h49;
mem[5323] = 8'h7d;
mem[5324] = 8'hcd;
mem[5325] = 8'h1c;
mem[5326] = 8'h02;
mem[5327] = 8'hd0;
mem[5328] = 8'hfe;
mem[5329] = 8'ha9;
mem[5330] = 8'hff;
mem[5331] = 8'h48;
mem[5332] = 8'h28;
mem[5333] = 8'ha4;
mem[5334] = 8'h14;
mem[5335] = 8'h08;
mem[5336] = 8'h98;
mem[5337] = 8'h49;
mem[5338] = 8'hc3;
mem[5339] = 8'ha8;
mem[5340] = 8'h28;
mem[5341] = 8'h8c;
mem[5342] = 8'h04;
mem[5343] = 8'h02;
mem[5344] = 8'h08;
mem[5345] = 8'h49;
mem[5346] = 8'hc3;
mem[5347] = 8'ha8;
mem[5348] = 8'hc0;
mem[5349] = 8'h82;
mem[5350] = 8'hd0;
mem[5351] = 8'hfe;
mem[5352] = 8'h68;
mem[5353] = 8'h09;
mem[5354] = 8'h08;
mem[5355] = 8'h49;
mem[5356] = 8'h7d;
mem[5357] = 8'hcd;
mem[5358] = 8'h1d;
mem[5359] = 8'h02;
mem[5360] = 8'hd0;
mem[5361] = 8'hfe;
mem[5362] = 8'ha9;
mem[5363] = 8'hff;
mem[5364] = 8'h48;
mem[5365] = 8'h28;
mem[5366] = 8'ha4;
mem[5367] = 8'h15;
mem[5368] = 8'h08;
mem[5369] = 8'h98;
mem[5370] = 8'h49;
mem[5371] = 8'hc3;
mem[5372] = 8'ha8;
mem[5373] = 8'h28;
mem[5374] = 8'h8c;
mem[5375] = 8'h05;
mem[5376] = 8'h02;
mem[5377] = 8'h08;
mem[5378] = 8'h49;
mem[5379] = 8'hc3;
mem[5380] = 8'ha8;
mem[5381] = 8'hc0;
mem[5382] = 8'h41;
mem[5383] = 8'hd0;
mem[5384] = 8'hfe;
mem[5385] = 8'h68;
mem[5386] = 8'h09;
mem[5387] = 8'h08;
mem[5388] = 8'h49;
mem[5389] = 8'h7d;
mem[5390] = 8'hcd;
mem[5391] = 8'h1e;
mem[5392] = 8'h02;
mem[5393] = 8'hd0;
mem[5394] = 8'hfe;
mem[5395] = 8'ha9;
mem[5396] = 8'hff;
mem[5397] = 8'h48;
mem[5398] = 8'h28;
mem[5399] = 8'ha4;
mem[5400] = 8'h16;
mem[5401] = 8'h08;
mem[5402] = 8'h98;
mem[5403] = 8'h49;
mem[5404] = 8'hc3;
mem[5405] = 8'ha8;
mem[5406] = 8'h28;
mem[5407] = 8'h8c;
mem[5408] = 8'h06;
mem[5409] = 8'h02;
mem[5410] = 8'h08;
mem[5411] = 8'h49;
mem[5412] = 8'hc3;
mem[5413] = 8'ha8;
mem[5414] = 8'hc0;
mem[5415] = 8'h00;
mem[5416] = 8'hd0;
mem[5417] = 8'hfe;
mem[5418] = 8'h68;
mem[5419] = 8'h09;
mem[5420] = 8'h08;
mem[5421] = 8'h49;
mem[5422] = 8'h7d;
mem[5423] = 8'hcd;
mem[5424] = 8'h1f;
mem[5425] = 8'h02;
mem[5426] = 8'hd0;
mem[5427] = 8'hfe;
mem[5428] = 8'ha9;
mem[5429] = 8'h00;
mem[5430] = 8'h48;
mem[5431] = 8'h28;
mem[5432] = 8'hac;
mem[5433] = 8'h17;
mem[5434] = 8'h02;
mem[5435] = 8'h08;
mem[5436] = 8'h98;
mem[5437] = 8'h49;
mem[5438] = 8'hc3;
mem[5439] = 8'ha8;
mem[5440] = 8'h28;
mem[5441] = 8'h84;
mem[5442] = 8'h0c;
mem[5443] = 8'h08;
mem[5444] = 8'h49;
mem[5445] = 8'hc3;
mem[5446] = 8'ha8;
mem[5447] = 8'hc4;
mem[5448] = 8'h13;
mem[5449] = 8'hd0;
mem[5450] = 8'hfe;
mem[5451] = 8'h68;
mem[5452] = 8'h09;
mem[5453] = 8'h08;
mem[5454] = 8'h49;
mem[5455] = 8'h38;
mem[5456] = 8'hcd;
mem[5457] = 8'h1c;
mem[5458] = 8'h02;
mem[5459] = 8'hd0;
mem[5460] = 8'hfe;
mem[5461] = 8'ha9;
mem[5462] = 8'h00;
mem[5463] = 8'h48;
mem[5464] = 8'h28;
mem[5465] = 8'hac;
mem[5466] = 8'h18;
mem[5467] = 8'h02;
mem[5468] = 8'h08;
mem[5469] = 8'h98;
mem[5470] = 8'h49;
mem[5471] = 8'hc3;
mem[5472] = 8'ha8;
mem[5473] = 8'h28;
mem[5474] = 8'h84;
mem[5475] = 8'h0d;
mem[5476] = 8'h08;
mem[5477] = 8'h49;
mem[5478] = 8'hc3;
mem[5479] = 8'ha8;
mem[5480] = 8'hc4;
mem[5481] = 8'h14;
mem[5482] = 8'hd0;
mem[5483] = 8'hfe;
mem[5484] = 8'h68;
mem[5485] = 8'h09;
mem[5486] = 8'h08;
mem[5487] = 8'h49;
mem[5488] = 8'h38;
mem[5489] = 8'hcd;
mem[5490] = 8'h1d;
mem[5491] = 8'h02;
mem[5492] = 8'hd0;
mem[5493] = 8'hfe;
mem[5494] = 8'ha9;
mem[5495] = 8'h00;
mem[5496] = 8'h48;
mem[5497] = 8'h28;
mem[5498] = 8'hac;
mem[5499] = 8'h19;
mem[5500] = 8'h02;
mem[5501] = 8'h08;
mem[5502] = 8'h98;
mem[5503] = 8'h49;
mem[5504] = 8'hc3;
mem[5505] = 8'ha8;
mem[5506] = 8'h28;
mem[5507] = 8'h84;
mem[5508] = 8'h0e;
mem[5509] = 8'h08;
mem[5510] = 8'h49;
mem[5511] = 8'hc3;
mem[5512] = 8'ha8;
mem[5513] = 8'hc4;
mem[5514] = 8'h15;
mem[5515] = 8'hd0;
mem[5516] = 8'hfe;
mem[5517] = 8'h68;
mem[5518] = 8'h09;
mem[5519] = 8'h08;
mem[5520] = 8'h49;
mem[5521] = 8'h38;
mem[5522] = 8'hcd;
mem[5523] = 8'h1e;
mem[5524] = 8'h02;
mem[5525] = 8'hd0;
mem[5526] = 8'hfe;
mem[5527] = 8'ha9;
mem[5528] = 8'h00;
mem[5529] = 8'h48;
mem[5530] = 8'h28;
mem[5531] = 8'hac;
mem[5532] = 8'h1a;
mem[5533] = 8'h02;
mem[5534] = 8'h08;
mem[5535] = 8'h98;
mem[5536] = 8'h49;
mem[5537] = 8'hc3;
mem[5538] = 8'ha8;
mem[5539] = 8'h28;
mem[5540] = 8'h84;
mem[5541] = 8'h0f;
mem[5542] = 8'h08;
mem[5543] = 8'h49;
mem[5544] = 8'hc3;
mem[5545] = 8'ha8;
mem[5546] = 8'hc4;
mem[5547] = 8'h16;
mem[5548] = 8'hd0;
mem[5549] = 8'hfe;
mem[5550] = 8'h68;
mem[5551] = 8'h09;
mem[5552] = 8'h08;
mem[5553] = 8'h49;
mem[5554] = 8'h38;
mem[5555] = 8'hcd;
mem[5556] = 8'h1f;
mem[5557] = 8'h02;
mem[5558] = 8'hd0;
mem[5559] = 8'hfe;
mem[5560] = 8'ha9;
mem[5561] = 8'hff;
mem[5562] = 8'h48;
mem[5563] = 8'h28;
mem[5564] = 8'hac;
mem[5565] = 8'h17;
mem[5566] = 8'h02;
mem[5567] = 8'h08;
mem[5568] = 8'h98;
mem[5569] = 8'h49;
mem[5570] = 8'hc3;
mem[5571] = 8'ha8;
mem[5572] = 8'h28;
mem[5573] = 8'h84;
mem[5574] = 8'h0c;
mem[5575] = 8'h08;
mem[5576] = 8'h49;
mem[5577] = 8'hc3;
mem[5578] = 8'ha8;
mem[5579] = 8'hc5;
mem[5580] = 8'h13;
mem[5581] = 8'hd0;
mem[5582] = 8'hfe;
mem[5583] = 8'h68;
mem[5584] = 8'h09;
mem[5585] = 8'h08;
mem[5586] = 8'h49;
mem[5587] = 8'h7d;
mem[5588] = 8'hcd;
mem[5589] = 8'h1c;
mem[5590] = 8'h02;
mem[5591] = 8'hd0;
mem[5592] = 8'hfe;
mem[5593] = 8'ha9;
mem[5594] = 8'hff;
mem[5595] = 8'h48;
mem[5596] = 8'h28;
mem[5597] = 8'hac;
mem[5598] = 8'h18;
mem[5599] = 8'h02;
mem[5600] = 8'h08;
mem[5601] = 8'h98;
mem[5602] = 8'h49;
mem[5603] = 8'hc3;
mem[5604] = 8'ha8;
mem[5605] = 8'h28;
mem[5606] = 8'h84;
mem[5607] = 8'h0d;
mem[5608] = 8'h08;
mem[5609] = 8'h49;
mem[5610] = 8'hc3;
mem[5611] = 8'ha8;
mem[5612] = 8'hc5;
mem[5613] = 8'h14;
mem[5614] = 8'hd0;
mem[5615] = 8'hfe;
mem[5616] = 8'h68;
mem[5617] = 8'h09;
mem[5618] = 8'h08;
mem[5619] = 8'h49;
mem[5620] = 8'h7d;
mem[5621] = 8'hcd;
mem[5622] = 8'h1d;
mem[5623] = 8'h02;
mem[5624] = 8'hd0;
mem[5625] = 8'hfe;
mem[5626] = 8'ha9;
mem[5627] = 8'hff;
mem[5628] = 8'h48;
mem[5629] = 8'h28;
mem[5630] = 8'hac;
mem[5631] = 8'h19;
mem[5632] = 8'h02;
mem[5633] = 8'h08;
mem[5634] = 8'h98;
mem[5635] = 8'h49;
mem[5636] = 8'hc3;
mem[5637] = 8'ha8;
mem[5638] = 8'h28;
mem[5639] = 8'h84;
mem[5640] = 8'h0e;
mem[5641] = 8'h08;
mem[5642] = 8'h49;
mem[5643] = 8'hc3;
mem[5644] = 8'ha8;
mem[5645] = 8'hc5;
mem[5646] = 8'h15;
mem[5647] = 8'hd0;
mem[5648] = 8'hfe;
mem[5649] = 8'h68;
mem[5650] = 8'h09;
mem[5651] = 8'h08;
mem[5652] = 8'h49;
mem[5653] = 8'h7d;
mem[5654] = 8'hcd;
mem[5655] = 8'h1e;
mem[5656] = 8'h02;
mem[5657] = 8'hd0;
mem[5658] = 8'hfe;
mem[5659] = 8'ha9;
mem[5660] = 8'hff;
mem[5661] = 8'h48;
mem[5662] = 8'h28;
mem[5663] = 8'hac;
mem[5664] = 8'h1a;
mem[5665] = 8'h02;
mem[5666] = 8'h08;
mem[5667] = 8'h98;
mem[5668] = 8'h49;
mem[5669] = 8'hc3;
mem[5670] = 8'ha8;
mem[5671] = 8'h28;
mem[5672] = 8'h84;
mem[5673] = 8'h0f;
mem[5674] = 8'h08;
mem[5675] = 8'h49;
mem[5676] = 8'hc3;
mem[5677] = 8'ha8;
mem[5678] = 8'hc5;
mem[5679] = 8'h16;
mem[5680] = 8'hd0;
mem[5681] = 8'hfe;
mem[5682] = 8'h68;
mem[5683] = 8'h09;
mem[5684] = 8'h08;
mem[5685] = 8'h49;
mem[5686] = 8'h7d;
mem[5687] = 8'hcd;
mem[5688] = 8'h1f;
mem[5689] = 8'h02;
mem[5690] = 8'hd0;
mem[5691] = 8'hfe;
mem[5692] = 8'ha9;
mem[5693] = 8'h00;
mem[5694] = 8'h48;
mem[5695] = 8'h28;
mem[5696] = 8'ha0;
mem[5697] = 8'hc3;
mem[5698] = 8'h08;
mem[5699] = 8'hcc;
mem[5700] = 8'h17;
mem[5701] = 8'h02;
mem[5702] = 8'hd0;
mem[5703] = 8'hfe;
mem[5704] = 8'h68;
mem[5705] = 8'h09;
mem[5706] = 8'h08;
mem[5707] = 8'h49;
mem[5708] = 8'h38;
mem[5709] = 8'hcd;
mem[5710] = 8'h1c;
mem[5711] = 8'h02;
mem[5712] = 8'hd0;
mem[5713] = 8'hfe;
mem[5714] = 8'ha9;
mem[5715] = 8'h00;
mem[5716] = 8'h48;
mem[5717] = 8'h28;
mem[5718] = 8'ha0;
mem[5719] = 8'h82;
mem[5720] = 8'h08;
mem[5721] = 8'hcc;
mem[5722] = 8'h18;
mem[5723] = 8'h02;
mem[5724] = 8'hd0;
mem[5725] = 8'hfe;
mem[5726] = 8'h68;
mem[5727] = 8'h09;
mem[5728] = 8'h08;
mem[5729] = 8'h49;
mem[5730] = 8'h38;
mem[5731] = 8'hcd;
mem[5732] = 8'h1d;
mem[5733] = 8'h02;
mem[5734] = 8'hd0;
mem[5735] = 8'hfe;
mem[5736] = 8'ha9;
mem[5737] = 8'h00;
mem[5738] = 8'h48;
mem[5739] = 8'h28;
mem[5740] = 8'ha0;
mem[5741] = 8'h41;
mem[5742] = 8'h08;
mem[5743] = 8'hcc;
mem[5744] = 8'h19;
mem[5745] = 8'h02;
mem[5746] = 8'hd0;
mem[5747] = 8'hfe;
mem[5748] = 8'h68;
mem[5749] = 8'h09;
mem[5750] = 8'h08;
mem[5751] = 8'h49;
mem[5752] = 8'h38;
mem[5753] = 8'hcd;
mem[5754] = 8'h1e;
mem[5755] = 8'h02;
mem[5756] = 8'hd0;
mem[5757] = 8'hfe;
mem[5758] = 8'ha9;
mem[5759] = 8'h00;
mem[5760] = 8'h48;
mem[5761] = 8'h28;
mem[5762] = 8'ha0;
mem[5763] = 8'h00;
mem[5764] = 8'h08;
mem[5765] = 8'hcc;
mem[5766] = 8'h1a;
mem[5767] = 8'h02;
mem[5768] = 8'hd0;
mem[5769] = 8'hfe;
mem[5770] = 8'h68;
mem[5771] = 8'h09;
mem[5772] = 8'h08;
mem[5773] = 8'h49;
mem[5774] = 8'h38;
mem[5775] = 8'hcd;
mem[5776] = 8'h1f;
mem[5777] = 8'h02;
mem[5778] = 8'hd0;
mem[5779] = 8'hfe;
mem[5780] = 8'ha9;
mem[5781] = 8'hff;
mem[5782] = 8'h48;
mem[5783] = 8'h28;
mem[5784] = 8'ha0;
mem[5785] = 8'hc3;
mem[5786] = 8'h08;
mem[5787] = 8'hcc;
mem[5788] = 8'h17;
mem[5789] = 8'h02;
mem[5790] = 8'hd0;
mem[5791] = 8'hfe;
mem[5792] = 8'h68;
mem[5793] = 8'h09;
mem[5794] = 8'h08;
mem[5795] = 8'h49;
mem[5796] = 8'h7d;
mem[5797] = 8'hcd;
mem[5798] = 8'h1c;
mem[5799] = 8'h02;
mem[5800] = 8'hd0;
mem[5801] = 8'hfe;
mem[5802] = 8'ha9;
mem[5803] = 8'hff;
mem[5804] = 8'h48;
mem[5805] = 8'h28;
mem[5806] = 8'ha0;
mem[5807] = 8'h82;
mem[5808] = 8'h08;
mem[5809] = 8'hcc;
mem[5810] = 8'h18;
mem[5811] = 8'h02;
mem[5812] = 8'hd0;
mem[5813] = 8'hfe;
mem[5814] = 8'h68;
mem[5815] = 8'h09;
mem[5816] = 8'h08;
mem[5817] = 8'h49;
mem[5818] = 8'h7d;
mem[5819] = 8'hcd;
mem[5820] = 8'h1d;
mem[5821] = 8'h02;
mem[5822] = 8'hd0;
mem[5823] = 8'hfe;
mem[5824] = 8'ha9;
mem[5825] = 8'hff;
mem[5826] = 8'h48;
mem[5827] = 8'h28;
mem[5828] = 8'ha0;
mem[5829] = 8'h41;
mem[5830] = 8'h08;
mem[5831] = 8'hcc;
mem[5832] = 8'h19;
mem[5833] = 8'h02;
mem[5834] = 8'hd0;
mem[5835] = 8'hfe;
mem[5836] = 8'h68;
mem[5837] = 8'h09;
mem[5838] = 8'h08;
mem[5839] = 8'h49;
mem[5840] = 8'h7d;
mem[5841] = 8'hcd;
mem[5842] = 8'h1e;
mem[5843] = 8'h02;
mem[5844] = 8'hd0;
mem[5845] = 8'hfe;
mem[5846] = 8'ha9;
mem[5847] = 8'hff;
mem[5848] = 8'h48;
mem[5849] = 8'h28;
mem[5850] = 8'ha0;
mem[5851] = 8'h00;
mem[5852] = 8'h08;
mem[5853] = 8'hcc;
mem[5854] = 8'h1a;
mem[5855] = 8'h02;
mem[5856] = 8'hd0;
mem[5857] = 8'hfe;
mem[5858] = 8'h68;
mem[5859] = 8'h09;
mem[5860] = 8'h08;
mem[5861] = 8'h49;
mem[5862] = 8'h7d;
mem[5863] = 8'hcd;
mem[5864] = 8'h1f;
mem[5865] = 8'h02;
mem[5866] = 8'hd0;
mem[5867] = 8'hfe;
mem[5868] = 8'ha0;
mem[5869] = 8'h00;
mem[5870] = 8'ha5;
mem[5871] = 8'h0c;
mem[5872] = 8'h49;
mem[5873] = 8'hc3;
mem[5874] = 8'hc5;
mem[5875] = 8'h13;
mem[5876] = 8'hd0;
mem[5877] = 8'hfe;
mem[5878] = 8'h84;
mem[5879] = 8'h0c;
mem[5880] = 8'had;
mem[5881] = 8'h03;
mem[5882] = 8'h02;
mem[5883] = 8'h49;
mem[5884] = 8'hc3;
mem[5885] = 8'hcd;
mem[5886] = 8'h17;
mem[5887] = 8'h02;
mem[5888] = 8'hd0;
mem[5889] = 8'hfe;
mem[5890] = 8'h8c;
mem[5891] = 8'h03;
mem[5892] = 8'h02;
mem[5893] = 8'ha5;
mem[5894] = 8'h0d;
mem[5895] = 8'h49;
mem[5896] = 8'hc3;
mem[5897] = 8'hc5;
mem[5898] = 8'h14;
mem[5899] = 8'hd0;
mem[5900] = 8'hfe;
mem[5901] = 8'h84;
mem[5902] = 8'h0d;
mem[5903] = 8'had;
mem[5904] = 8'h04;
mem[5905] = 8'h02;
mem[5906] = 8'h49;
mem[5907] = 8'hc3;
mem[5908] = 8'hcd;
mem[5909] = 8'h18;
mem[5910] = 8'h02;
mem[5911] = 8'hd0;
mem[5912] = 8'hfe;
mem[5913] = 8'h8c;
mem[5914] = 8'h04;
mem[5915] = 8'h02;
mem[5916] = 8'ha5;
mem[5917] = 8'h0e;
mem[5918] = 8'h49;
mem[5919] = 8'hc3;
mem[5920] = 8'hc5;
mem[5921] = 8'h15;
mem[5922] = 8'hd0;
mem[5923] = 8'hfe;
mem[5924] = 8'h84;
mem[5925] = 8'h0e;
mem[5926] = 8'had;
mem[5927] = 8'h05;
mem[5928] = 8'h02;
mem[5929] = 8'h49;
mem[5930] = 8'hc3;
mem[5931] = 8'hcd;
mem[5932] = 8'h19;
mem[5933] = 8'h02;
mem[5934] = 8'hd0;
mem[5935] = 8'hfe;
mem[5936] = 8'h8c;
mem[5937] = 8'h05;
mem[5938] = 8'h02;
mem[5939] = 8'ha5;
mem[5940] = 8'h0f;
mem[5941] = 8'h49;
mem[5942] = 8'hc3;
mem[5943] = 8'hc5;
mem[5944] = 8'h16;
mem[5945] = 8'hd0;
mem[5946] = 8'hfe;
mem[5947] = 8'h84;
mem[5948] = 8'h0f;
mem[5949] = 8'had;
mem[5950] = 8'h06;
mem[5951] = 8'h02;
mem[5952] = 8'h49;
mem[5953] = 8'hc3;
mem[5954] = 8'hcd;
mem[5955] = 8'h1a;
mem[5956] = 8'h02;
mem[5957] = 8'hd0;
mem[5958] = 8'hfe;
mem[5959] = 8'h8c;
mem[5960] = 8'h06;
mem[5961] = 8'h02;
mem[5962] = 8'had;
mem[5963] = 8'h00;
mem[5964] = 8'h02;
mem[5965] = 8'hc9;
mem[5966] = 8'h14;
mem[5967] = 8'hd0;
mem[5968] = 8'hfe;
mem[5969] = 8'ha9;
mem[5970] = 8'h15;
mem[5971] = 8'h8d;
mem[5972] = 8'h00;
mem[5973] = 8'h02;
mem[5974] = 8'ha2;
mem[5975] = 8'h03;
mem[5976] = 8'ha9;
mem[5977] = 8'h00;
mem[5978] = 8'h48;
mem[5979] = 8'h28;
mem[5980] = 8'hb5;
mem[5981] = 8'h13;
mem[5982] = 8'h08;
mem[5983] = 8'h49;
mem[5984] = 8'hc3;
mem[5985] = 8'h28;
mem[5986] = 8'h9d;
mem[5987] = 8'h03;
mem[5988] = 8'h02;
mem[5989] = 8'h08;
mem[5990] = 8'h49;
mem[5991] = 8'hc3;
mem[5992] = 8'hdd;
mem[5993] = 8'h17;
mem[5994] = 8'h02;
mem[5995] = 8'hd0;
mem[5996] = 8'hfe;
mem[5997] = 8'h68;
mem[5998] = 8'h09;
mem[5999] = 8'h08;
mem[6000] = 8'h49;
mem[6001] = 8'h38;
mem[6002] = 8'hdd;
mem[6003] = 8'h1c;
mem[6004] = 8'h02;
mem[6005] = 8'hd0;
mem[6006] = 8'hfe;
mem[6007] = 8'hca;
mem[6008] = 8'h10;
mem[6009] = 8'hde;
mem[6010] = 8'ha2;
mem[6011] = 8'h03;
mem[6012] = 8'ha9;
mem[6013] = 8'hff;
mem[6014] = 8'h48;
mem[6015] = 8'h28;
mem[6016] = 8'hb5;
mem[6017] = 8'h13;
mem[6018] = 8'h08;
mem[6019] = 8'h49;
mem[6020] = 8'hc3;
mem[6021] = 8'h28;
mem[6022] = 8'h9d;
mem[6023] = 8'h03;
mem[6024] = 8'h02;
mem[6025] = 8'h08;
mem[6026] = 8'h49;
mem[6027] = 8'hc3;
mem[6028] = 8'hdd;
mem[6029] = 8'h17;
mem[6030] = 8'h02;
mem[6031] = 8'hd0;
mem[6032] = 8'hfe;
mem[6033] = 8'h68;
mem[6034] = 8'h09;
mem[6035] = 8'h08;
mem[6036] = 8'h49;
mem[6037] = 8'h7d;
mem[6038] = 8'hdd;
mem[6039] = 8'h1c;
mem[6040] = 8'h02;
mem[6041] = 8'hd0;
mem[6042] = 8'hfe;
mem[6043] = 8'hca;
mem[6044] = 8'h10;
mem[6045] = 8'hde;
mem[6046] = 8'ha2;
mem[6047] = 8'h03;
mem[6048] = 8'ha9;
mem[6049] = 8'h00;
mem[6050] = 8'h48;
mem[6051] = 8'h28;
mem[6052] = 8'hbd;
mem[6053] = 8'h17;
mem[6054] = 8'h02;
mem[6055] = 8'h08;
mem[6056] = 8'h49;
mem[6057] = 8'hc3;
mem[6058] = 8'h28;
mem[6059] = 8'h95;
mem[6060] = 8'h0c;
mem[6061] = 8'h08;
mem[6062] = 8'h49;
mem[6063] = 8'hc3;
mem[6064] = 8'hd5;
mem[6065] = 8'h13;
mem[6066] = 8'hd0;
mem[6067] = 8'hfe;
mem[6068] = 8'h68;
mem[6069] = 8'h09;
mem[6070] = 8'h08;
mem[6071] = 8'h49;
mem[6072] = 8'h38;
mem[6073] = 8'hdd;
mem[6074] = 8'h1c;
mem[6075] = 8'h02;
mem[6076] = 8'hd0;
mem[6077] = 8'hfe;
mem[6078] = 8'hca;
mem[6079] = 8'h10;
mem[6080] = 8'hdf;
mem[6081] = 8'ha2;
mem[6082] = 8'h03;
mem[6083] = 8'ha9;
mem[6084] = 8'hff;
mem[6085] = 8'h48;
mem[6086] = 8'h28;
mem[6087] = 8'hbd;
mem[6088] = 8'h17;
mem[6089] = 8'h02;
mem[6090] = 8'h08;
mem[6091] = 8'h49;
mem[6092] = 8'hc3;
mem[6093] = 8'h28;
mem[6094] = 8'h95;
mem[6095] = 8'h0c;
mem[6096] = 8'h08;
mem[6097] = 8'h49;
mem[6098] = 8'hc3;
mem[6099] = 8'hd5;
mem[6100] = 8'h13;
mem[6101] = 8'hd0;
mem[6102] = 8'hfe;
mem[6103] = 8'h68;
mem[6104] = 8'h09;
mem[6105] = 8'h08;
mem[6106] = 8'h49;
mem[6107] = 8'h7d;
mem[6108] = 8'hdd;
mem[6109] = 8'h1c;
mem[6110] = 8'h02;
mem[6111] = 8'hd0;
mem[6112] = 8'hfe;
mem[6113] = 8'hca;
mem[6114] = 8'h10;
mem[6115] = 8'hdf;
mem[6116] = 8'ha2;
mem[6117] = 8'h03;
mem[6118] = 8'ha0;
mem[6119] = 8'h00;
mem[6120] = 8'hb5;
mem[6121] = 8'h0c;
mem[6122] = 8'h49;
mem[6123] = 8'hc3;
mem[6124] = 8'hd5;
mem[6125] = 8'h13;
mem[6126] = 8'hd0;
mem[6127] = 8'hfe;
mem[6128] = 8'h94;
mem[6129] = 8'h0c;
mem[6130] = 8'hbd;
mem[6131] = 8'h03;
mem[6132] = 8'h02;
mem[6133] = 8'h49;
mem[6134] = 8'hc3;
mem[6135] = 8'hdd;
mem[6136] = 8'h17;
mem[6137] = 8'h02;
mem[6138] = 8'hd0;
mem[6139] = 8'hfe;
mem[6140] = 8'h8a;
mem[6141] = 8'h9d;
mem[6142] = 8'h03;
mem[6143] = 8'h02;
mem[6144] = 8'hca;
mem[6145] = 8'h10;
mem[6146] = 8'he5;
mem[6147] = 8'had;
mem[6148] = 8'h00;
mem[6149] = 8'h02;
mem[6150] = 8'hc9;
mem[6151] = 8'h15;
mem[6152] = 8'hd0;
mem[6153] = 8'hfe;
mem[6154] = 8'ha9;
mem[6155] = 8'h16;
mem[6156] = 8'h8d;
mem[6157] = 8'h00;
mem[6158] = 8'h02;
mem[6159] = 8'ha0;
mem[6160] = 8'h03;
mem[6161] = 8'ha9;
mem[6162] = 8'h00;
mem[6163] = 8'h48;
mem[6164] = 8'h28;
mem[6165] = 8'hb1;
mem[6166] = 8'h24;
mem[6167] = 8'h08;
mem[6168] = 8'h49;
mem[6169] = 8'hc3;
mem[6170] = 8'h28;
mem[6171] = 8'h99;
mem[6172] = 8'h03;
mem[6173] = 8'h02;
mem[6174] = 8'h08;
mem[6175] = 8'h49;
mem[6176] = 8'hc3;
mem[6177] = 8'hd9;
mem[6178] = 8'h17;
mem[6179] = 8'h02;
mem[6180] = 8'hd0;
mem[6181] = 8'hfe;
mem[6182] = 8'h68;
mem[6183] = 8'h09;
mem[6184] = 8'h08;
mem[6185] = 8'h49;
mem[6186] = 8'h38;
mem[6187] = 8'hd9;
mem[6188] = 8'h1c;
mem[6189] = 8'h02;
mem[6190] = 8'hd0;
mem[6191] = 8'hfe;
mem[6192] = 8'h88;
mem[6193] = 8'h10;
mem[6194] = 8'hde;
mem[6195] = 8'ha0;
mem[6196] = 8'h03;
mem[6197] = 8'ha9;
mem[6198] = 8'hff;
mem[6199] = 8'h48;
mem[6200] = 8'h28;
mem[6201] = 8'hb1;
mem[6202] = 8'h24;
mem[6203] = 8'h08;
mem[6204] = 8'h49;
mem[6205] = 8'hc3;
mem[6206] = 8'h28;
mem[6207] = 8'h99;
mem[6208] = 8'h03;
mem[6209] = 8'h02;
mem[6210] = 8'h08;
mem[6211] = 8'h49;
mem[6212] = 8'hc3;
mem[6213] = 8'hd9;
mem[6214] = 8'h17;
mem[6215] = 8'h02;
mem[6216] = 8'hd0;
mem[6217] = 8'hfe;
mem[6218] = 8'h68;
mem[6219] = 8'h09;
mem[6220] = 8'h08;
mem[6221] = 8'h49;
mem[6222] = 8'h7d;
mem[6223] = 8'hd9;
mem[6224] = 8'h1c;
mem[6225] = 8'h02;
mem[6226] = 8'hd0;
mem[6227] = 8'hfe;
mem[6228] = 8'h88;
mem[6229] = 8'h10;
mem[6230] = 8'hde;
mem[6231] = 8'ha0;
mem[6232] = 8'h03;
mem[6233] = 8'ha2;
mem[6234] = 8'h00;
mem[6235] = 8'hb9;
mem[6236] = 8'h03;
mem[6237] = 8'h02;
mem[6238] = 8'h49;
mem[6239] = 8'hc3;
mem[6240] = 8'hd9;
mem[6241] = 8'h17;
mem[6242] = 8'h02;
mem[6243] = 8'hd0;
mem[6244] = 8'hfe;
mem[6245] = 8'h8a;
mem[6246] = 8'h99;
mem[6247] = 8'h03;
mem[6248] = 8'h02;
mem[6249] = 8'h88;
mem[6250] = 8'h10;
mem[6251] = 8'hef;
mem[6252] = 8'ha0;
mem[6253] = 8'h03;
mem[6254] = 8'ha9;
mem[6255] = 8'h00;
mem[6256] = 8'h48;
mem[6257] = 8'h28;
mem[6258] = 8'hb9;
mem[6259] = 8'h17;
mem[6260] = 8'h02;
mem[6261] = 8'h08;
mem[6262] = 8'h49;
mem[6263] = 8'hc3;
mem[6264] = 8'h28;
mem[6265] = 8'h91;
mem[6266] = 8'h30;
mem[6267] = 8'h08;
mem[6268] = 8'h49;
mem[6269] = 8'hc3;
mem[6270] = 8'hd1;
mem[6271] = 8'h24;
mem[6272] = 8'hd0;
mem[6273] = 8'hfe;
mem[6274] = 8'h68;
mem[6275] = 8'h09;
mem[6276] = 8'h08;
mem[6277] = 8'h49;
mem[6278] = 8'h38;
mem[6279] = 8'hd9;
mem[6280] = 8'h1c;
mem[6281] = 8'h02;
mem[6282] = 8'hd0;
mem[6283] = 8'hfe;
mem[6284] = 8'h88;
mem[6285] = 8'h10;
mem[6286] = 8'hdf;
mem[6287] = 8'ha0;
mem[6288] = 8'h03;
mem[6289] = 8'ha9;
mem[6290] = 8'hff;
mem[6291] = 8'h48;
mem[6292] = 8'h28;
mem[6293] = 8'hb9;
mem[6294] = 8'h17;
mem[6295] = 8'h02;
mem[6296] = 8'h08;
mem[6297] = 8'h49;
mem[6298] = 8'hc3;
mem[6299] = 8'h28;
mem[6300] = 8'h91;
mem[6301] = 8'h30;
mem[6302] = 8'h08;
mem[6303] = 8'h49;
mem[6304] = 8'hc3;
mem[6305] = 8'hd1;
mem[6306] = 8'h24;
mem[6307] = 8'hd0;
mem[6308] = 8'hfe;
mem[6309] = 8'h68;
mem[6310] = 8'h09;
mem[6311] = 8'h08;
mem[6312] = 8'h49;
mem[6313] = 8'h7d;
mem[6314] = 8'hd9;
mem[6315] = 8'h1c;
mem[6316] = 8'h02;
mem[6317] = 8'hd0;
mem[6318] = 8'hfe;
mem[6319] = 8'h88;
mem[6320] = 8'h10;
mem[6321] = 8'hdf;
mem[6322] = 8'ha0;
mem[6323] = 8'h03;
mem[6324] = 8'ha2;
mem[6325] = 8'h00;
mem[6326] = 8'hb9;
mem[6327] = 8'h03;
mem[6328] = 8'h02;
mem[6329] = 8'h49;
mem[6330] = 8'hc3;
mem[6331] = 8'hd9;
mem[6332] = 8'h17;
mem[6333] = 8'h02;
mem[6334] = 8'hd0;
mem[6335] = 8'hfe;
mem[6336] = 8'h8a;
mem[6337] = 8'h99;
mem[6338] = 8'h03;
mem[6339] = 8'h02;
mem[6340] = 8'h88;
mem[6341] = 8'h10;
mem[6342] = 8'hef;
mem[6343] = 8'ha2;
mem[6344] = 8'h06;
mem[6345] = 8'ha0;
mem[6346] = 8'h03;
mem[6347] = 8'ha9;
mem[6348] = 8'h00;
mem[6349] = 8'h48;
mem[6350] = 8'h28;
mem[6351] = 8'ha1;
mem[6352] = 8'h24;
mem[6353] = 8'h08;
mem[6354] = 8'h49;
mem[6355] = 8'hc3;
mem[6356] = 8'h28;
mem[6357] = 8'h81;
mem[6358] = 8'h30;
mem[6359] = 8'h08;
mem[6360] = 8'h49;
mem[6361] = 8'hc3;
mem[6362] = 8'hd9;
mem[6363] = 8'h17;
mem[6364] = 8'h02;
mem[6365] = 8'hd0;
mem[6366] = 8'hfe;
mem[6367] = 8'h68;
mem[6368] = 8'h09;
mem[6369] = 8'h08;
mem[6370] = 8'h49;
mem[6371] = 8'h38;
mem[6372] = 8'hd9;
mem[6373] = 8'h1c;
mem[6374] = 8'h02;
mem[6375] = 8'hd0;
mem[6376] = 8'hfe;
mem[6377] = 8'hca;
mem[6378] = 8'hca;
mem[6379] = 8'h88;
mem[6380] = 8'h10;
mem[6381] = 8'hdd;
mem[6382] = 8'ha2;
mem[6383] = 8'h06;
mem[6384] = 8'ha0;
mem[6385] = 8'h03;
mem[6386] = 8'ha9;
mem[6387] = 8'hff;
mem[6388] = 8'h48;
mem[6389] = 8'h28;
mem[6390] = 8'ha1;
mem[6391] = 8'h24;
mem[6392] = 8'h08;
mem[6393] = 8'h49;
mem[6394] = 8'hc3;
mem[6395] = 8'h28;
mem[6396] = 8'h81;
mem[6397] = 8'h30;
mem[6398] = 8'h08;
mem[6399] = 8'h49;
mem[6400] = 8'hc3;
mem[6401] = 8'hd9;
mem[6402] = 8'h17;
mem[6403] = 8'h02;
mem[6404] = 8'hd0;
mem[6405] = 8'hfe;
mem[6406] = 8'h68;
mem[6407] = 8'h09;
mem[6408] = 8'h08;
mem[6409] = 8'h49;
mem[6410] = 8'h7d;
mem[6411] = 8'hd9;
mem[6412] = 8'h1c;
mem[6413] = 8'h02;
mem[6414] = 8'hd0;
mem[6415] = 8'hfe;
mem[6416] = 8'hca;
mem[6417] = 8'hca;
mem[6418] = 8'h88;
mem[6419] = 8'h10;
mem[6420] = 8'hdd;
mem[6421] = 8'ha0;
mem[6422] = 8'h03;
mem[6423] = 8'ha2;
mem[6424] = 8'h00;
mem[6425] = 8'hb9;
mem[6426] = 8'h03;
mem[6427] = 8'h02;
mem[6428] = 8'h49;
mem[6429] = 8'hc3;
mem[6430] = 8'hd9;
mem[6431] = 8'h17;
mem[6432] = 8'h02;
mem[6433] = 8'hd0;
mem[6434] = 8'hfe;
mem[6435] = 8'h8a;
mem[6436] = 8'h99;
mem[6437] = 8'h03;
mem[6438] = 8'h02;
mem[6439] = 8'h88;
mem[6440] = 8'h10;
mem[6441] = 8'hef;
mem[6442] = 8'had;
mem[6443] = 8'h00;
mem[6444] = 8'h02;
mem[6445] = 8'hc9;
mem[6446] = 8'h16;
mem[6447] = 8'hd0;
mem[6448] = 8'hfe;
mem[6449] = 8'ha9;
mem[6450] = 8'h17;
mem[6451] = 8'h8d;
mem[6452] = 8'h00;
mem[6453] = 8'h02;
mem[6454] = 8'ha2;
mem[6455] = 8'hfd;
mem[6456] = 8'hb5;
mem[6457] = 8'h19;
mem[6458] = 8'h9d;
mem[6459] = 8'h09;
mem[6460] = 8'h01;
mem[6461] = 8'hca;
mem[6462] = 8'he0;
mem[6463] = 8'hfa;
mem[6464] = 8'hb0;
mem[6465] = 8'hf6;
mem[6466] = 8'ha2;
mem[6467] = 8'hfd;
mem[6468] = 8'hbd;
mem[6469] = 8'h1d;
mem[6470] = 8'h01;
mem[6471] = 8'h95;
mem[6472] = 8'h12;
mem[6473] = 8'hca;
mem[6474] = 8'he0;
mem[6475] = 8'hfa;
mem[6476] = 8'hb0;
mem[6477] = 8'hf6;
mem[6478] = 8'ha2;
mem[6479] = 8'h03;
mem[6480] = 8'ha0;
mem[6481] = 8'h00;
mem[6482] = 8'hb5;
mem[6483] = 8'h0c;
mem[6484] = 8'hd5;
mem[6485] = 8'h13;
mem[6486] = 8'hd0;
mem[6487] = 8'hfe;
mem[6488] = 8'h94;
mem[6489] = 8'h0c;
mem[6490] = 8'hbd;
mem[6491] = 8'h03;
mem[6492] = 8'h02;
mem[6493] = 8'hdd;
mem[6494] = 8'h17;
mem[6495] = 8'h02;
mem[6496] = 8'hd0;
mem[6497] = 8'hfe;
mem[6498] = 8'h8a;
mem[6499] = 8'h9d;
mem[6500] = 8'h03;
mem[6501] = 8'h02;
mem[6502] = 8'hca;
mem[6503] = 8'h10;
mem[6504] = 8'he9;
mem[6505] = 8'ha0;
mem[6506] = 8'hfb;
mem[6507] = 8'ha2;
mem[6508] = 8'hfe;
mem[6509] = 8'ha1;
mem[6510] = 8'h2c;
mem[6511] = 8'h99;
mem[6512] = 8'h0b;
mem[6513] = 8'h01;
mem[6514] = 8'hca;
mem[6515] = 8'hca;
mem[6516] = 8'h88;
mem[6517] = 8'hc0;
mem[6518] = 8'hf8;
mem[6519] = 8'hb0;
mem[6520] = 8'hf4;
mem[6521] = 8'ha0;
mem[6522] = 8'h03;
mem[6523] = 8'ha2;
mem[6524] = 8'h00;
mem[6525] = 8'hb9;
mem[6526] = 8'h03;
mem[6527] = 8'h02;
mem[6528] = 8'hd9;
mem[6529] = 8'h17;
mem[6530] = 8'h02;
mem[6531] = 8'hd0;
mem[6532] = 8'hfe;
mem[6533] = 8'h8a;
mem[6534] = 8'h99;
mem[6535] = 8'h03;
mem[6536] = 8'h02;
mem[6537] = 8'h88;
mem[6538] = 8'h10;
mem[6539] = 8'hf1;
mem[6540] = 8'ha0;
mem[6541] = 8'hfb;
mem[6542] = 8'hb9;
mem[6543] = 8'h1f;
mem[6544] = 8'h01;
mem[6545] = 8'h91;
mem[6546] = 8'h38;
mem[6547] = 8'h88;
mem[6548] = 8'hc0;
mem[6549] = 8'hf8;
mem[6550] = 8'hb0;
mem[6551] = 8'hf6;
mem[6552] = 8'ha0;
mem[6553] = 8'h03;
mem[6554] = 8'ha2;
mem[6555] = 8'h00;
mem[6556] = 8'hb9;
mem[6557] = 8'h03;
mem[6558] = 8'h02;
mem[6559] = 8'hd9;
mem[6560] = 8'h17;
mem[6561] = 8'h02;
mem[6562] = 8'hd0;
mem[6563] = 8'hfe;
mem[6564] = 8'h8a;
mem[6565] = 8'h99;
mem[6566] = 8'h03;
mem[6567] = 8'h02;
mem[6568] = 8'h88;
mem[6569] = 8'h10;
mem[6570] = 8'hf1;
mem[6571] = 8'ha0;
mem[6572] = 8'hfb;
mem[6573] = 8'ha2;
mem[6574] = 8'hfe;
mem[6575] = 8'hb1;
mem[6576] = 8'h2e;
mem[6577] = 8'h81;
mem[6578] = 8'h38;
mem[6579] = 8'hca;
mem[6580] = 8'hca;
mem[6581] = 8'h88;
mem[6582] = 8'hc0;
mem[6583] = 8'hf8;
mem[6584] = 8'hb0;
mem[6585] = 8'hf5;
mem[6586] = 8'ha0;
mem[6587] = 8'h03;
mem[6588] = 8'ha2;
mem[6589] = 8'h00;
mem[6590] = 8'hb9;
mem[6591] = 8'h03;
mem[6592] = 8'h02;
mem[6593] = 8'hd9;
mem[6594] = 8'h17;
mem[6595] = 8'h02;
mem[6596] = 8'hd0;
mem[6597] = 8'hfe;
mem[6598] = 8'h8a;
mem[6599] = 8'h99;
mem[6600] = 8'h03;
mem[6601] = 8'h02;
mem[6602] = 8'h88;
mem[6603] = 8'h10;
mem[6604] = 8'hf1;
mem[6605] = 8'had;
mem[6606] = 8'h00;
mem[6607] = 8'h02;
mem[6608] = 8'hc9;
mem[6609] = 8'h17;
mem[6610] = 8'hd0;
mem[6611] = 8'hfe;
mem[6612] = 8'ha9;
mem[6613] = 8'h18;
mem[6614] = 8'h8d;
mem[6615] = 8'h00;
mem[6616] = 8'h02;
mem[6617] = 8'ha9;
mem[6618] = 8'h00;
mem[6619] = 8'h48;
mem[6620] = 8'h28;
mem[6621] = 8'ha5;
mem[6622] = 8'h13;
mem[6623] = 8'h08;
mem[6624] = 8'h49;
mem[6625] = 8'hc3;
mem[6626] = 8'h28;
mem[6627] = 8'h8d;
mem[6628] = 8'h03;
mem[6629] = 8'h02;
mem[6630] = 8'h08;
mem[6631] = 8'h49;
mem[6632] = 8'hc3;
mem[6633] = 8'hc9;
mem[6634] = 8'hc3;
mem[6635] = 8'hd0;
mem[6636] = 8'hfe;
mem[6637] = 8'h68;
mem[6638] = 8'h09;
mem[6639] = 8'h08;
mem[6640] = 8'h49;
mem[6641] = 8'h38;
mem[6642] = 8'hcd;
mem[6643] = 8'h1c;
mem[6644] = 8'h02;
mem[6645] = 8'hd0;
mem[6646] = 8'hfe;
mem[6647] = 8'ha9;
mem[6648] = 8'h00;
mem[6649] = 8'h48;
mem[6650] = 8'h28;
mem[6651] = 8'ha5;
mem[6652] = 8'h14;
mem[6653] = 8'h08;
mem[6654] = 8'h49;
mem[6655] = 8'hc3;
mem[6656] = 8'h28;
mem[6657] = 8'h8d;
mem[6658] = 8'h04;
mem[6659] = 8'h02;
mem[6660] = 8'h08;
mem[6661] = 8'h49;
mem[6662] = 8'hc3;
mem[6663] = 8'hc9;
mem[6664] = 8'h82;
mem[6665] = 8'hd0;
mem[6666] = 8'hfe;
mem[6667] = 8'h68;
mem[6668] = 8'h09;
mem[6669] = 8'h08;
mem[6670] = 8'h49;
mem[6671] = 8'h38;
mem[6672] = 8'hcd;
mem[6673] = 8'h1d;
mem[6674] = 8'h02;
mem[6675] = 8'hd0;
mem[6676] = 8'hfe;
mem[6677] = 8'ha9;
mem[6678] = 8'h00;
mem[6679] = 8'h48;
mem[6680] = 8'h28;
mem[6681] = 8'ha5;
mem[6682] = 8'h15;
mem[6683] = 8'h08;
mem[6684] = 8'h49;
mem[6685] = 8'hc3;
mem[6686] = 8'h28;
mem[6687] = 8'h8d;
mem[6688] = 8'h05;
mem[6689] = 8'h02;
mem[6690] = 8'h08;
mem[6691] = 8'h49;
mem[6692] = 8'hc3;
mem[6693] = 8'hc9;
mem[6694] = 8'h41;
mem[6695] = 8'hd0;
mem[6696] = 8'hfe;
mem[6697] = 8'h68;
mem[6698] = 8'h09;
mem[6699] = 8'h08;
mem[6700] = 8'h49;
mem[6701] = 8'h38;
mem[6702] = 8'hcd;
mem[6703] = 8'h1e;
mem[6704] = 8'h02;
mem[6705] = 8'hd0;
mem[6706] = 8'hfe;
mem[6707] = 8'ha9;
mem[6708] = 8'h00;
mem[6709] = 8'h48;
mem[6710] = 8'h28;
mem[6711] = 8'ha5;
mem[6712] = 8'h16;
mem[6713] = 8'h08;
mem[6714] = 8'h49;
mem[6715] = 8'hc3;
mem[6716] = 8'h28;
mem[6717] = 8'h8d;
mem[6718] = 8'h06;
mem[6719] = 8'h02;
mem[6720] = 8'h08;
mem[6721] = 8'h49;
mem[6722] = 8'hc3;
mem[6723] = 8'hc9;
mem[6724] = 8'h00;
mem[6725] = 8'hd0;
mem[6726] = 8'hfe;
mem[6727] = 8'h68;
mem[6728] = 8'h09;
mem[6729] = 8'h08;
mem[6730] = 8'h49;
mem[6731] = 8'h38;
mem[6732] = 8'hcd;
mem[6733] = 8'h1f;
mem[6734] = 8'h02;
mem[6735] = 8'hd0;
mem[6736] = 8'hfe;
mem[6737] = 8'ha9;
mem[6738] = 8'hff;
mem[6739] = 8'h48;
mem[6740] = 8'h28;
mem[6741] = 8'ha5;
mem[6742] = 8'h13;
mem[6743] = 8'h08;
mem[6744] = 8'h49;
mem[6745] = 8'hc3;
mem[6746] = 8'h28;
mem[6747] = 8'h8d;
mem[6748] = 8'h03;
mem[6749] = 8'h02;
mem[6750] = 8'h08;
mem[6751] = 8'h49;
mem[6752] = 8'hc3;
mem[6753] = 8'hc9;
mem[6754] = 8'hc3;
mem[6755] = 8'hd0;
mem[6756] = 8'hfe;
mem[6757] = 8'h68;
mem[6758] = 8'h09;
mem[6759] = 8'h08;
mem[6760] = 8'h49;
mem[6761] = 8'h7d;
mem[6762] = 8'hcd;
mem[6763] = 8'h1c;
mem[6764] = 8'h02;
mem[6765] = 8'hd0;
mem[6766] = 8'hfe;
mem[6767] = 8'ha9;
mem[6768] = 8'hff;
mem[6769] = 8'h48;
mem[6770] = 8'h28;
mem[6771] = 8'ha5;
mem[6772] = 8'h14;
mem[6773] = 8'h08;
mem[6774] = 8'h49;
mem[6775] = 8'hc3;
mem[6776] = 8'h28;
mem[6777] = 8'h8d;
mem[6778] = 8'h04;
mem[6779] = 8'h02;
mem[6780] = 8'h08;
mem[6781] = 8'h49;
mem[6782] = 8'hc3;
mem[6783] = 8'hc9;
mem[6784] = 8'h82;
mem[6785] = 8'hd0;
mem[6786] = 8'hfe;
mem[6787] = 8'h68;
mem[6788] = 8'h09;
mem[6789] = 8'h08;
mem[6790] = 8'h49;
mem[6791] = 8'h7d;
mem[6792] = 8'hcd;
mem[6793] = 8'h1d;
mem[6794] = 8'h02;
mem[6795] = 8'hd0;
mem[6796] = 8'hfe;
mem[6797] = 8'ha9;
mem[6798] = 8'hff;
mem[6799] = 8'h48;
mem[6800] = 8'h28;
mem[6801] = 8'ha5;
mem[6802] = 8'h15;
mem[6803] = 8'h08;
mem[6804] = 8'h49;
mem[6805] = 8'hc3;
mem[6806] = 8'h28;
mem[6807] = 8'h8d;
mem[6808] = 8'h05;
mem[6809] = 8'h02;
mem[6810] = 8'h08;
mem[6811] = 8'h49;
mem[6812] = 8'hc3;
mem[6813] = 8'hc9;
mem[6814] = 8'h41;
mem[6815] = 8'hd0;
mem[6816] = 8'hfe;
mem[6817] = 8'h68;
mem[6818] = 8'h09;
mem[6819] = 8'h08;
mem[6820] = 8'h49;
mem[6821] = 8'h7d;
mem[6822] = 8'hcd;
mem[6823] = 8'h1e;
mem[6824] = 8'h02;
mem[6825] = 8'hd0;
mem[6826] = 8'hfe;
mem[6827] = 8'ha9;
mem[6828] = 8'hff;
mem[6829] = 8'h48;
mem[6830] = 8'h28;
mem[6831] = 8'ha5;
mem[6832] = 8'h16;
mem[6833] = 8'h08;
mem[6834] = 8'h49;
mem[6835] = 8'hc3;
mem[6836] = 8'h28;
mem[6837] = 8'h8d;
mem[6838] = 8'h06;
mem[6839] = 8'h02;
mem[6840] = 8'h08;
mem[6841] = 8'h49;
mem[6842] = 8'hc3;
mem[6843] = 8'hc9;
mem[6844] = 8'h00;
mem[6845] = 8'hd0;
mem[6846] = 8'hfe;
mem[6847] = 8'h68;
mem[6848] = 8'h09;
mem[6849] = 8'h08;
mem[6850] = 8'h49;
mem[6851] = 8'h7d;
mem[6852] = 8'hcd;
mem[6853] = 8'h1f;
mem[6854] = 8'h02;
mem[6855] = 8'hd0;
mem[6856] = 8'hfe;
mem[6857] = 8'ha9;
mem[6858] = 8'h00;
mem[6859] = 8'h48;
mem[6860] = 8'h28;
mem[6861] = 8'had;
mem[6862] = 8'h17;
mem[6863] = 8'h02;
mem[6864] = 8'h08;
mem[6865] = 8'h49;
mem[6866] = 8'hc3;
mem[6867] = 8'h28;
mem[6868] = 8'h85;
mem[6869] = 8'h0c;
mem[6870] = 8'h08;
mem[6871] = 8'h49;
mem[6872] = 8'hc3;
mem[6873] = 8'hc5;
mem[6874] = 8'h13;
mem[6875] = 8'hd0;
mem[6876] = 8'hfe;
mem[6877] = 8'h68;
mem[6878] = 8'h09;
mem[6879] = 8'h08;
mem[6880] = 8'h49;
mem[6881] = 8'h38;
mem[6882] = 8'hcd;
mem[6883] = 8'h1c;
mem[6884] = 8'h02;
mem[6885] = 8'hd0;
mem[6886] = 8'hfe;
mem[6887] = 8'ha9;
mem[6888] = 8'h00;
mem[6889] = 8'h48;
mem[6890] = 8'h28;
mem[6891] = 8'had;
mem[6892] = 8'h18;
mem[6893] = 8'h02;
mem[6894] = 8'h08;
mem[6895] = 8'h49;
mem[6896] = 8'hc3;
mem[6897] = 8'h28;
mem[6898] = 8'h85;
mem[6899] = 8'h0d;
mem[6900] = 8'h08;
mem[6901] = 8'h49;
mem[6902] = 8'hc3;
mem[6903] = 8'hc5;
mem[6904] = 8'h14;
mem[6905] = 8'hd0;
mem[6906] = 8'hfe;
mem[6907] = 8'h68;
mem[6908] = 8'h09;
mem[6909] = 8'h08;
mem[6910] = 8'h49;
mem[6911] = 8'h38;
mem[6912] = 8'hcd;
mem[6913] = 8'h1d;
mem[6914] = 8'h02;
mem[6915] = 8'hd0;
mem[6916] = 8'hfe;
mem[6917] = 8'ha9;
mem[6918] = 8'h00;
mem[6919] = 8'h48;
mem[6920] = 8'h28;
mem[6921] = 8'had;
mem[6922] = 8'h19;
mem[6923] = 8'h02;
mem[6924] = 8'h08;
mem[6925] = 8'h49;
mem[6926] = 8'hc3;
mem[6927] = 8'h28;
mem[6928] = 8'h85;
mem[6929] = 8'h0e;
mem[6930] = 8'h08;
mem[6931] = 8'h49;
mem[6932] = 8'hc3;
mem[6933] = 8'hc5;
mem[6934] = 8'h15;
mem[6935] = 8'hd0;
mem[6936] = 8'hfe;
mem[6937] = 8'h68;
mem[6938] = 8'h09;
mem[6939] = 8'h08;
mem[6940] = 8'h49;
mem[6941] = 8'h38;
mem[6942] = 8'hcd;
mem[6943] = 8'h1e;
mem[6944] = 8'h02;
mem[6945] = 8'hd0;
mem[6946] = 8'hfe;
mem[6947] = 8'ha9;
mem[6948] = 8'h00;
mem[6949] = 8'h48;
mem[6950] = 8'h28;
mem[6951] = 8'had;
mem[6952] = 8'h1a;
mem[6953] = 8'h02;
mem[6954] = 8'h08;
mem[6955] = 8'h49;
mem[6956] = 8'hc3;
mem[6957] = 8'h28;
mem[6958] = 8'h85;
mem[6959] = 8'h0f;
mem[6960] = 8'h08;
mem[6961] = 8'h49;
mem[6962] = 8'hc3;
mem[6963] = 8'hc5;
mem[6964] = 8'h16;
mem[6965] = 8'hd0;
mem[6966] = 8'hfe;
mem[6967] = 8'h68;
mem[6968] = 8'h09;
mem[6969] = 8'h08;
mem[6970] = 8'h49;
mem[6971] = 8'h38;
mem[6972] = 8'hcd;
mem[6973] = 8'h1f;
mem[6974] = 8'h02;
mem[6975] = 8'hd0;
mem[6976] = 8'hfe;
mem[6977] = 8'ha9;
mem[6978] = 8'hff;
mem[6979] = 8'h48;
mem[6980] = 8'h28;
mem[6981] = 8'had;
mem[6982] = 8'h17;
mem[6983] = 8'h02;
mem[6984] = 8'h08;
mem[6985] = 8'h49;
mem[6986] = 8'hc3;
mem[6987] = 8'h28;
mem[6988] = 8'h85;
mem[6989] = 8'h0c;
mem[6990] = 8'h08;
mem[6991] = 8'h49;
mem[6992] = 8'hc3;
mem[6993] = 8'hc5;
mem[6994] = 8'h13;
mem[6995] = 8'hd0;
mem[6996] = 8'hfe;
mem[6997] = 8'h68;
mem[6998] = 8'h09;
mem[6999] = 8'h08;
mem[7000] = 8'h49;
mem[7001] = 8'h7d;
mem[7002] = 8'hcd;
mem[7003] = 8'h1c;
mem[7004] = 8'h02;
mem[7005] = 8'hd0;
mem[7006] = 8'hfe;
mem[7007] = 8'ha9;
mem[7008] = 8'hff;
mem[7009] = 8'h48;
mem[7010] = 8'h28;
mem[7011] = 8'had;
mem[7012] = 8'h18;
mem[7013] = 8'h02;
mem[7014] = 8'h08;
mem[7015] = 8'h49;
mem[7016] = 8'hc3;
mem[7017] = 8'h28;
mem[7018] = 8'h85;
mem[7019] = 8'h0d;
mem[7020] = 8'h08;
mem[7021] = 8'h49;
mem[7022] = 8'hc3;
mem[7023] = 8'hc5;
mem[7024] = 8'h14;
mem[7025] = 8'hd0;
mem[7026] = 8'hfe;
mem[7027] = 8'h68;
mem[7028] = 8'h09;
mem[7029] = 8'h08;
mem[7030] = 8'h49;
mem[7031] = 8'h7d;
mem[7032] = 8'hcd;
mem[7033] = 8'h1d;
mem[7034] = 8'h02;
mem[7035] = 8'hd0;
mem[7036] = 8'hfe;
mem[7037] = 8'ha9;
mem[7038] = 8'hff;
mem[7039] = 8'h48;
mem[7040] = 8'h28;
mem[7041] = 8'had;
mem[7042] = 8'h19;
mem[7043] = 8'h02;
mem[7044] = 8'h08;
mem[7045] = 8'h49;
mem[7046] = 8'hc3;
mem[7047] = 8'h28;
mem[7048] = 8'h85;
mem[7049] = 8'h0e;
mem[7050] = 8'h08;
mem[7051] = 8'h49;
mem[7052] = 8'hc3;
mem[7053] = 8'hc5;
mem[7054] = 8'h15;
mem[7055] = 8'hd0;
mem[7056] = 8'hfe;
mem[7057] = 8'h68;
mem[7058] = 8'h09;
mem[7059] = 8'h08;
mem[7060] = 8'h49;
mem[7061] = 8'h7d;
mem[7062] = 8'hcd;
mem[7063] = 8'h1e;
mem[7064] = 8'h02;
mem[7065] = 8'hd0;
mem[7066] = 8'hfe;
mem[7067] = 8'ha9;
mem[7068] = 8'hff;
mem[7069] = 8'h48;
mem[7070] = 8'h28;
mem[7071] = 8'had;
mem[7072] = 8'h1a;
mem[7073] = 8'h02;
mem[7074] = 8'h08;
mem[7075] = 8'h49;
mem[7076] = 8'hc3;
mem[7077] = 8'h28;
mem[7078] = 8'h85;
mem[7079] = 8'h0f;
mem[7080] = 8'h08;
mem[7081] = 8'h49;
mem[7082] = 8'hc3;
mem[7083] = 8'hc5;
mem[7084] = 8'h16;
mem[7085] = 8'hd0;
mem[7086] = 8'hfe;
mem[7087] = 8'h68;
mem[7088] = 8'h09;
mem[7089] = 8'h08;
mem[7090] = 8'h49;
mem[7091] = 8'h7d;
mem[7092] = 8'hcd;
mem[7093] = 8'h1f;
mem[7094] = 8'h02;
mem[7095] = 8'hd0;
mem[7096] = 8'hfe;
mem[7097] = 8'ha9;
mem[7098] = 8'h00;
mem[7099] = 8'h48;
mem[7100] = 8'h28;
mem[7101] = 8'ha9;
mem[7102] = 8'hc3;
mem[7103] = 8'h08;
mem[7104] = 8'hcd;
mem[7105] = 8'h17;
mem[7106] = 8'h02;
mem[7107] = 8'hd0;
mem[7108] = 8'hfe;
mem[7109] = 8'h68;
mem[7110] = 8'h09;
mem[7111] = 8'h08;
mem[7112] = 8'h49;
mem[7113] = 8'h38;
mem[7114] = 8'hcd;
mem[7115] = 8'h1c;
mem[7116] = 8'h02;
mem[7117] = 8'hd0;
mem[7118] = 8'hfe;
mem[7119] = 8'ha9;
mem[7120] = 8'h00;
mem[7121] = 8'h48;
mem[7122] = 8'h28;
mem[7123] = 8'ha9;
mem[7124] = 8'h82;
mem[7125] = 8'h08;
mem[7126] = 8'hcd;
mem[7127] = 8'h18;
mem[7128] = 8'h02;
mem[7129] = 8'hd0;
mem[7130] = 8'hfe;
mem[7131] = 8'h68;
mem[7132] = 8'h09;
mem[7133] = 8'h08;
mem[7134] = 8'h49;
mem[7135] = 8'h38;
mem[7136] = 8'hcd;
mem[7137] = 8'h1d;
mem[7138] = 8'h02;
mem[7139] = 8'hd0;
mem[7140] = 8'hfe;
mem[7141] = 8'ha9;
mem[7142] = 8'h00;
mem[7143] = 8'h48;
mem[7144] = 8'h28;
mem[7145] = 8'ha9;
mem[7146] = 8'h41;
mem[7147] = 8'h08;
mem[7148] = 8'hcd;
mem[7149] = 8'h19;
mem[7150] = 8'h02;
mem[7151] = 8'hd0;
mem[7152] = 8'hfe;
mem[7153] = 8'h68;
mem[7154] = 8'h09;
mem[7155] = 8'h08;
mem[7156] = 8'h49;
mem[7157] = 8'h38;
mem[7158] = 8'hcd;
mem[7159] = 8'h1e;
mem[7160] = 8'h02;
mem[7161] = 8'hd0;
mem[7162] = 8'hfe;
mem[7163] = 8'ha9;
mem[7164] = 8'h00;
mem[7165] = 8'h48;
mem[7166] = 8'h28;
mem[7167] = 8'ha9;
mem[7168] = 8'h00;
mem[7169] = 8'h08;
mem[7170] = 8'hcd;
mem[7171] = 8'h1a;
mem[7172] = 8'h02;
mem[7173] = 8'hd0;
mem[7174] = 8'hfe;
mem[7175] = 8'h68;
mem[7176] = 8'h09;
mem[7177] = 8'h08;
mem[7178] = 8'h49;
mem[7179] = 8'h38;
mem[7180] = 8'hcd;
mem[7181] = 8'h1f;
mem[7182] = 8'h02;
mem[7183] = 8'hd0;
mem[7184] = 8'hfe;
mem[7185] = 8'ha9;
mem[7186] = 8'hff;
mem[7187] = 8'h48;
mem[7188] = 8'h28;
mem[7189] = 8'ha9;
mem[7190] = 8'hc3;
mem[7191] = 8'h08;
mem[7192] = 8'hcd;
mem[7193] = 8'h17;
mem[7194] = 8'h02;
mem[7195] = 8'hd0;
mem[7196] = 8'hfe;
mem[7197] = 8'h68;
mem[7198] = 8'h09;
mem[7199] = 8'h08;
mem[7200] = 8'h49;
mem[7201] = 8'h7d;
mem[7202] = 8'hcd;
mem[7203] = 8'h1c;
mem[7204] = 8'h02;
mem[7205] = 8'hd0;
mem[7206] = 8'hfe;
mem[7207] = 8'ha9;
mem[7208] = 8'hff;
mem[7209] = 8'h48;
mem[7210] = 8'h28;
mem[7211] = 8'ha9;
mem[7212] = 8'h82;
mem[7213] = 8'h08;
mem[7214] = 8'hcd;
mem[7215] = 8'h18;
mem[7216] = 8'h02;
mem[7217] = 8'hd0;
mem[7218] = 8'hfe;
mem[7219] = 8'h68;
mem[7220] = 8'h09;
mem[7221] = 8'h08;
mem[7222] = 8'h49;
mem[7223] = 8'h7d;
mem[7224] = 8'hcd;
mem[7225] = 8'h1d;
mem[7226] = 8'h02;
mem[7227] = 8'hd0;
mem[7228] = 8'hfe;
mem[7229] = 8'ha9;
mem[7230] = 8'hff;
mem[7231] = 8'h48;
mem[7232] = 8'h28;
mem[7233] = 8'ha9;
mem[7234] = 8'h41;
mem[7235] = 8'h08;
mem[7236] = 8'hcd;
mem[7237] = 8'h19;
mem[7238] = 8'h02;
mem[7239] = 8'hd0;
mem[7240] = 8'hfe;
mem[7241] = 8'h68;
mem[7242] = 8'h09;
mem[7243] = 8'h08;
mem[7244] = 8'h49;
mem[7245] = 8'h7d;
mem[7246] = 8'hcd;
mem[7247] = 8'h1e;
mem[7248] = 8'h02;
mem[7249] = 8'hd0;
mem[7250] = 8'hfe;
mem[7251] = 8'ha9;
mem[7252] = 8'hff;
mem[7253] = 8'h48;
mem[7254] = 8'h28;
mem[7255] = 8'ha9;
mem[7256] = 8'h00;
mem[7257] = 8'h08;
mem[7258] = 8'hcd;
mem[7259] = 8'h1a;
mem[7260] = 8'h02;
mem[7261] = 8'hd0;
mem[7262] = 8'hfe;
mem[7263] = 8'h68;
mem[7264] = 8'h09;
mem[7265] = 8'h08;
mem[7266] = 8'h49;
mem[7267] = 8'h7d;
mem[7268] = 8'hcd;
mem[7269] = 8'h1f;
mem[7270] = 8'h02;
mem[7271] = 8'hd0;
mem[7272] = 8'hfe;
mem[7273] = 8'ha2;
mem[7274] = 8'h00;
mem[7275] = 8'ha5;
mem[7276] = 8'h0c;
mem[7277] = 8'h49;
mem[7278] = 8'hc3;
mem[7279] = 8'hc5;
mem[7280] = 8'h13;
mem[7281] = 8'hd0;
mem[7282] = 8'hfe;
mem[7283] = 8'h86;
mem[7284] = 8'h0c;
mem[7285] = 8'had;
mem[7286] = 8'h03;
mem[7287] = 8'h02;
mem[7288] = 8'h49;
mem[7289] = 8'hc3;
mem[7290] = 8'hcd;
mem[7291] = 8'h17;
mem[7292] = 8'h02;
mem[7293] = 8'hd0;
mem[7294] = 8'hfe;
mem[7295] = 8'h8e;
mem[7296] = 8'h03;
mem[7297] = 8'h02;
mem[7298] = 8'ha5;
mem[7299] = 8'h0d;
mem[7300] = 8'h49;
mem[7301] = 8'hc3;
mem[7302] = 8'hc5;
mem[7303] = 8'h14;
mem[7304] = 8'hd0;
mem[7305] = 8'hfe;
mem[7306] = 8'h86;
mem[7307] = 8'h0d;
mem[7308] = 8'had;
mem[7309] = 8'h04;
mem[7310] = 8'h02;
mem[7311] = 8'h49;
mem[7312] = 8'hc3;
mem[7313] = 8'hcd;
mem[7314] = 8'h18;
mem[7315] = 8'h02;
mem[7316] = 8'hd0;
mem[7317] = 8'hfe;
mem[7318] = 8'h8e;
mem[7319] = 8'h04;
mem[7320] = 8'h02;
mem[7321] = 8'ha5;
mem[7322] = 8'h0e;
mem[7323] = 8'h49;
mem[7324] = 8'hc3;
mem[7325] = 8'hc5;
mem[7326] = 8'h15;
mem[7327] = 8'hd0;
mem[7328] = 8'hfe;
mem[7329] = 8'h86;
mem[7330] = 8'h0e;
mem[7331] = 8'had;
mem[7332] = 8'h05;
mem[7333] = 8'h02;
mem[7334] = 8'h49;
mem[7335] = 8'hc3;
mem[7336] = 8'hcd;
mem[7337] = 8'h19;
mem[7338] = 8'h02;
mem[7339] = 8'hd0;
mem[7340] = 8'hfe;
mem[7341] = 8'h8e;
mem[7342] = 8'h05;
mem[7343] = 8'h02;
mem[7344] = 8'ha5;
mem[7345] = 8'h0f;
mem[7346] = 8'h49;
mem[7347] = 8'hc3;
mem[7348] = 8'hc5;
mem[7349] = 8'h16;
mem[7350] = 8'hd0;
mem[7351] = 8'hfe;
mem[7352] = 8'h86;
mem[7353] = 8'h0f;
mem[7354] = 8'had;
mem[7355] = 8'h06;
mem[7356] = 8'h02;
mem[7357] = 8'h49;
mem[7358] = 8'hc3;
mem[7359] = 8'hcd;
mem[7360] = 8'h1a;
mem[7361] = 8'h02;
mem[7362] = 8'hd0;
mem[7363] = 8'hfe;
mem[7364] = 8'h8e;
mem[7365] = 8'h06;
mem[7366] = 8'h02;
mem[7367] = 8'had;
mem[7368] = 8'h00;
mem[7369] = 8'h02;
mem[7370] = 8'hc9;
mem[7371] = 8'h18;
mem[7372] = 8'hd0;
mem[7373] = 8'hfe;
mem[7374] = 8'ha9;
mem[7375] = 8'h19;
mem[7376] = 8'h8d;
mem[7377] = 8'h00;
mem[7378] = 8'h02;
mem[7379] = 8'ha9;
mem[7380] = 8'h00;
mem[7381] = 8'h48;
mem[7382] = 8'ha9;
mem[7383] = 8'hff;
mem[7384] = 8'h28;
mem[7385] = 8'h24;
mem[7386] = 8'h16;
mem[7387] = 8'h08;
mem[7388] = 8'hc9;
mem[7389] = 8'hff;
mem[7390] = 8'hd0;
mem[7391] = 8'hfe;
mem[7392] = 8'h68;
mem[7393] = 8'h48;
mem[7394] = 8'h09;
mem[7395] = 8'h08;
mem[7396] = 8'hc9;
mem[7397] = 8'h3a;
mem[7398] = 8'hd0;
mem[7399] = 8'hfe;
mem[7400] = 8'h28;
mem[7401] = 8'ha9;
mem[7402] = 8'h00;
mem[7403] = 8'h48;
mem[7404] = 8'ha9;
mem[7405] = 8'h01;
mem[7406] = 8'h28;
mem[7407] = 8'h24;
mem[7408] = 8'h15;
mem[7409] = 8'h08;
mem[7410] = 8'hc9;
mem[7411] = 8'h01;
mem[7412] = 8'hd0;
mem[7413] = 8'hfe;
mem[7414] = 8'h68;
mem[7415] = 8'h48;
mem[7416] = 8'h09;
mem[7417] = 8'h08;
mem[7418] = 8'hc9;
mem[7419] = 8'h78;
mem[7420] = 8'hd0;
mem[7421] = 8'hfe;
mem[7422] = 8'h28;
mem[7423] = 8'ha9;
mem[7424] = 8'h00;
mem[7425] = 8'h48;
mem[7426] = 8'ha9;
mem[7427] = 8'h01;
mem[7428] = 8'h28;
mem[7429] = 8'h24;
mem[7430] = 8'h14;
mem[7431] = 8'h08;
mem[7432] = 8'hc9;
mem[7433] = 8'h01;
mem[7434] = 8'hd0;
mem[7435] = 8'hfe;
mem[7436] = 8'h68;
mem[7437] = 8'h48;
mem[7438] = 8'h09;
mem[7439] = 8'h08;
mem[7440] = 8'hc9;
mem[7441] = 8'hba;
mem[7442] = 8'hd0;
mem[7443] = 8'hfe;
mem[7444] = 8'h28;
mem[7445] = 8'ha9;
mem[7446] = 8'h00;
mem[7447] = 8'h48;
mem[7448] = 8'ha9;
mem[7449] = 8'h01;
mem[7450] = 8'h28;
mem[7451] = 8'h24;
mem[7452] = 8'h13;
mem[7453] = 8'h08;
mem[7454] = 8'hc9;
mem[7455] = 8'h01;
mem[7456] = 8'hd0;
mem[7457] = 8'hfe;
mem[7458] = 8'h68;
mem[7459] = 8'h48;
mem[7460] = 8'h09;
mem[7461] = 8'h08;
mem[7462] = 8'hc9;
mem[7463] = 8'hf8;
mem[7464] = 8'hd0;
mem[7465] = 8'hfe;
mem[7466] = 8'h28;
mem[7467] = 8'ha9;
mem[7468] = 8'hff;
mem[7469] = 8'h48;
mem[7470] = 8'ha9;
mem[7471] = 8'hff;
mem[7472] = 8'h28;
mem[7473] = 8'h24;
mem[7474] = 8'h16;
mem[7475] = 8'h08;
mem[7476] = 8'hc9;
mem[7477] = 8'hff;
mem[7478] = 8'hd0;
mem[7479] = 8'hfe;
mem[7480] = 8'h68;
mem[7481] = 8'h48;
mem[7482] = 8'h09;
mem[7483] = 8'h08;
mem[7484] = 8'hc9;
mem[7485] = 8'h3f;
mem[7486] = 8'hd0;
mem[7487] = 8'hfe;
mem[7488] = 8'h28;
mem[7489] = 8'ha9;
mem[7490] = 8'hff;
mem[7491] = 8'h48;
mem[7492] = 8'ha9;
mem[7493] = 8'h01;
mem[7494] = 8'h28;
mem[7495] = 8'h24;
mem[7496] = 8'h15;
mem[7497] = 8'h08;
mem[7498] = 8'hc9;
mem[7499] = 8'h01;
mem[7500] = 8'hd0;
mem[7501] = 8'hfe;
mem[7502] = 8'h68;
mem[7503] = 8'h48;
mem[7504] = 8'h09;
mem[7505] = 8'h08;
mem[7506] = 8'hc9;
mem[7507] = 8'h7d;
mem[7508] = 8'hd0;
mem[7509] = 8'hfe;
mem[7510] = 8'h28;
mem[7511] = 8'ha9;
mem[7512] = 8'hff;
mem[7513] = 8'h48;
mem[7514] = 8'ha9;
mem[7515] = 8'h01;
mem[7516] = 8'h28;
mem[7517] = 8'h24;
mem[7518] = 8'h14;
mem[7519] = 8'h08;
mem[7520] = 8'hc9;
mem[7521] = 8'h01;
mem[7522] = 8'hd0;
mem[7523] = 8'hfe;
mem[7524] = 8'h68;
mem[7525] = 8'h48;
mem[7526] = 8'h09;
mem[7527] = 8'h08;
mem[7528] = 8'hc9;
mem[7529] = 8'hbf;
mem[7530] = 8'hd0;
mem[7531] = 8'hfe;
mem[7532] = 8'h28;
mem[7533] = 8'ha9;
mem[7534] = 8'hff;
mem[7535] = 8'h48;
mem[7536] = 8'ha9;
mem[7537] = 8'h01;
mem[7538] = 8'h28;
mem[7539] = 8'h24;
mem[7540] = 8'h13;
mem[7541] = 8'h08;
mem[7542] = 8'hc9;
mem[7543] = 8'h01;
mem[7544] = 8'hd0;
mem[7545] = 8'hfe;
mem[7546] = 8'h68;
mem[7547] = 8'h48;
mem[7548] = 8'h09;
mem[7549] = 8'h08;
mem[7550] = 8'hc9;
mem[7551] = 8'hfd;
mem[7552] = 8'hd0;
mem[7553] = 8'hfe;
mem[7554] = 8'h28;
mem[7555] = 8'ha9;
mem[7556] = 8'h00;
mem[7557] = 8'h48;
mem[7558] = 8'ha9;
mem[7559] = 8'hff;
mem[7560] = 8'h28;
mem[7561] = 8'h2c;
mem[7562] = 8'h1a;
mem[7563] = 8'h02;
mem[7564] = 8'h08;
mem[7565] = 8'hc9;
mem[7566] = 8'hff;
mem[7567] = 8'hd0;
mem[7568] = 8'hfe;
mem[7569] = 8'h68;
mem[7570] = 8'h48;
mem[7571] = 8'h09;
mem[7572] = 8'h08;
mem[7573] = 8'hc9;
mem[7574] = 8'h3a;
mem[7575] = 8'hd0;
mem[7576] = 8'hfe;
mem[7577] = 8'h28;
mem[7578] = 8'ha9;
mem[7579] = 8'h00;
mem[7580] = 8'h48;
mem[7581] = 8'ha9;
mem[7582] = 8'h01;
mem[7583] = 8'h28;
mem[7584] = 8'h2c;
mem[7585] = 8'h19;
mem[7586] = 8'h02;
mem[7587] = 8'h08;
mem[7588] = 8'hc9;
mem[7589] = 8'h01;
mem[7590] = 8'hd0;
mem[7591] = 8'hfe;
mem[7592] = 8'h68;
mem[7593] = 8'h48;
mem[7594] = 8'h09;
mem[7595] = 8'h08;
mem[7596] = 8'hc9;
mem[7597] = 8'h78;
mem[7598] = 8'hd0;
mem[7599] = 8'hfe;
mem[7600] = 8'h28;
mem[7601] = 8'ha9;
mem[7602] = 8'h00;
mem[7603] = 8'h48;
mem[7604] = 8'ha9;
mem[7605] = 8'h01;
mem[7606] = 8'h28;
mem[7607] = 8'h2c;
mem[7608] = 8'h18;
mem[7609] = 8'h02;
mem[7610] = 8'h08;
mem[7611] = 8'hc9;
mem[7612] = 8'h01;
mem[7613] = 8'hd0;
mem[7614] = 8'hfe;
mem[7615] = 8'h68;
mem[7616] = 8'h48;
mem[7617] = 8'h09;
mem[7618] = 8'h08;
mem[7619] = 8'hc9;
mem[7620] = 8'hba;
mem[7621] = 8'hd0;
mem[7622] = 8'hfe;
mem[7623] = 8'h28;
mem[7624] = 8'ha9;
mem[7625] = 8'h00;
mem[7626] = 8'h48;
mem[7627] = 8'ha9;
mem[7628] = 8'h01;
mem[7629] = 8'h28;
mem[7630] = 8'h2c;
mem[7631] = 8'h17;
mem[7632] = 8'h02;
mem[7633] = 8'h08;
mem[7634] = 8'hc9;
mem[7635] = 8'h01;
mem[7636] = 8'hd0;
mem[7637] = 8'hfe;
mem[7638] = 8'h68;
mem[7639] = 8'h48;
mem[7640] = 8'h09;
mem[7641] = 8'h08;
mem[7642] = 8'hc9;
mem[7643] = 8'hf8;
mem[7644] = 8'hd0;
mem[7645] = 8'hfe;
mem[7646] = 8'h28;
mem[7647] = 8'ha9;
mem[7648] = 8'hff;
mem[7649] = 8'h48;
mem[7650] = 8'ha9;
mem[7651] = 8'hff;
mem[7652] = 8'h28;
mem[7653] = 8'h2c;
mem[7654] = 8'h1a;
mem[7655] = 8'h02;
mem[7656] = 8'h08;
mem[7657] = 8'hc9;
mem[7658] = 8'hff;
mem[7659] = 8'hd0;
mem[7660] = 8'hfe;
mem[7661] = 8'h68;
mem[7662] = 8'h48;
mem[7663] = 8'h09;
mem[7664] = 8'h08;
mem[7665] = 8'hc9;
mem[7666] = 8'h3f;
mem[7667] = 8'hd0;
mem[7668] = 8'hfe;
mem[7669] = 8'h28;
mem[7670] = 8'ha9;
mem[7671] = 8'hff;
mem[7672] = 8'h48;
mem[7673] = 8'ha9;
mem[7674] = 8'h01;
mem[7675] = 8'h28;
mem[7676] = 8'h2c;
mem[7677] = 8'h19;
mem[7678] = 8'h02;
mem[7679] = 8'h08;
mem[7680] = 8'hc9;
mem[7681] = 8'h01;
mem[7682] = 8'hd0;
mem[7683] = 8'hfe;
mem[7684] = 8'h68;
mem[7685] = 8'h48;
mem[7686] = 8'h09;
mem[7687] = 8'h08;
mem[7688] = 8'hc9;
mem[7689] = 8'h7d;
mem[7690] = 8'hd0;
mem[7691] = 8'hfe;
mem[7692] = 8'h28;
mem[7693] = 8'ha9;
mem[7694] = 8'hff;
mem[7695] = 8'h48;
mem[7696] = 8'ha9;
mem[7697] = 8'h01;
mem[7698] = 8'h28;
mem[7699] = 8'h2c;
mem[7700] = 8'h18;
mem[7701] = 8'h02;
mem[7702] = 8'h08;
mem[7703] = 8'hc9;
mem[7704] = 8'h01;
mem[7705] = 8'hd0;
mem[7706] = 8'hfe;
mem[7707] = 8'h68;
mem[7708] = 8'h48;
mem[7709] = 8'h09;
mem[7710] = 8'h08;
mem[7711] = 8'hc9;
mem[7712] = 8'hbf;
mem[7713] = 8'hd0;
mem[7714] = 8'hfe;
mem[7715] = 8'h28;
mem[7716] = 8'ha9;
mem[7717] = 8'hff;
mem[7718] = 8'h48;
mem[7719] = 8'ha9;
mem[7720] = 8'h01;
mem[7721] = 8'h28;
mem[7722] = 8'h2c;
mem[7723] = 8'h17;
mem[7724] = 8'h02;
mem[7725] = 8'h08;
mem[7726] = 8'hc9;
mem[7727] = 8'h01;
mem[7728] = 8'hd0;
mem[7729] = 8'hfe;
mem[7730] = 8'h68;
mem[7731] = 8'h48;
mem[7732] = 8'h09;
mem[7733] = 8'h08;
mem[7734] = 8'hc9;
mem[7735] = 8'hfd;
mem[7736] = 8'hd0;
mem[7737] = 8'hfe;
mem[7738] = 8'h28;
mem[7739] = 8'had;
mem[7740] = 8'h00;
mem[7741] = 8'h02;
mem[7742] = 8'hc9;
mem[7743] = 8'h19;
mem[7744] = 8'hd0;
mem[7745] = 8'hfe;
mem[7746] = 8'ha9;
mem[7747] = 8'h1a;
mem[7748] = 8'h8d;
mem[7749] = 8'h00;
mem[7750] = 8'h02;
mem[7751] = 8'ha9;
mem[7752] = 8'h00;
mem[7753] = 8'h48;
mem[7754] = 8'ha2;
mem[7755] = 8'h80;
mem[7756] = 8'h28;
mem[7757] = 8'he4;
mem[7758] = 8'h17;
mem[7759] = 8'h08;
mem[7760] = 8'h68;
mem[7761] = 8'h48;
mem[7762] = 8'h09;
mem[7763] = 8'h08;
mem[7764] = 8'hc9;
mem[7765] = 8'h39;
mem[7766] = 8'hd0;
mem[7767] = 8'hfe;
mem[7768] = 8'h28;
mem[7769] = 8'hca;
mem[7770] = 8'he4;
mem[7771] = 8'h17;
mem[7772] = 8'h08;
mem[7773] = 8'h68;
mem[7774] = 8'h48;
mem[7775] = 8'h09;
mem[7776] = 8'h08;
mem[7777] = 8'hc9;
mem[7778] = 8'h3b;
mem[7779] = 8'hd0;
mem[7780] = 8'hfe;
mem[7781] = 8'h28;
mem[7782] = 8'hca;
mem[7783] = 8'he4;
mem[7784] = 8'h17;
mem[7785] = 8'h08;
mem[7786] = 8'he0;
mem[7787] = 8'h7e;
mem[7788] = 8'hd0;
mem[7789] = 8'hfe;
mem[7790] = 8'h68;
mem[7791] = 8'h48;
mem[7792] = 8'h09;
mem[7793] = 8'h08;
mem[7794] = 8'hc9;
mem[7795] = 8'hb8;
mem[7796] = 8'hd0;
mem[7797] = 8'hfe;
mem[7798] = 8'h28;
mem[7799] = 8'ha9;
mem[7800] = 8'hff;
mem[7801] = 8'h48;
mem[7802] = 8'ha2;
mem[7803] = 8'h80;
mem[7804] = 8'h28;
mem[7805] = 8'he4;
mem[7806] = 8'h17;
mem[7807] = 8'h08;
mem[7808] = 8'h68;
mem[7809] = 8'h48;
mem[7810] = 8'h09;
mem[7811] = 8'h08;
mem[7812] = 8'hc9;
mem[7813] = 8'h7d;
mem[7814] = 8'hd0;
mem[7815] = 8'hfe;
mem[7816] = 8'h28;
mem[7817] = 8'hca;
mem[7818] = 8'he4;
mem[7819] = 8'h17;
mem[7820] = 8'h08;
mem[7821] = 8'h68;
mem[7822] = 8'h48;
mem[7823] = 8'h09;
mem[7824] = 8'h08;
mem[7825] = 8'hc9;
mem[7826] = 8'h7f;
mem[7827] = 8'hd0;
mem[7828] = 8'hfe;
mem[7829] = 8'h28;
mem[7830] = 8'hca;
mem[7831] = 8'he4;
mem[7832] = 8'h17;
mem[7833] = 8'h08;
mem[7834] = 8'he0;
mem[7835] = 8'h7e;
mem[7836] = 8'hd0;
mem[7837] = 8'hfe;
mem[7838] = 8'h68;
mem[7839] = 8'h48;
mem[7840] = 8'h09;
mem[7841] = 8'h08;
mem[7842] = 8'hc9;
mem[7843] = 8'hfc;
mem[7844] = 8'hd0;
mem[7845] = 8'hfe;
mem[7846] = 8'h28;
mem[7847] = 8'ha9;
mem[7848] = 8'h00;
mem[7849] = 8'h48;
mem[7850] = 8'ha2;
mem[7851] = 8'h80;
mem[7852] = 8'h28;
mem[7853] = 8'hec;
mem[7854] = 8'h1b;
mem[7855] = 8'h02;
mem[7856] = 8'h08;
mem[7857] = 8'h68;
mem[7858] = 8'h48;
mem[7859] = 8'h09;
mem[7860] = 8'h08;
mem[7861] = 8'hc9;
mem[7862] = 8'h39;
mem[7863] = 8'hd0;
mem[7864] = 8'hfe;
mem[7865] = 8'h28;
mem[7866] = 8'hca;
mem[7867] = 8'hec;
mem[7868] = 8'h1b;
mem[7869] = 8'h02;
mem[7870] = 8'h08;
mem[7871] = 8'h68;
mem[7872] = 8'h48;
mem[7873] = 8'h09;
mem[7874] = 8'h08;
mem[7875] = 8'hc9;
mem[7876] = 8'h3b;
mem[7877] = 8'hd0;
mem[7878] = 8'hfe;
mem[7879] = 8'h28;
mem[7880] = 8'hca;
mem[7881] = 8'hec;
mem[7882] = 8'h1b;
mem[7883] = 8'h02;
mem[7884] = 8'h08;
mem[7885] = 8'he0;
mem[7886] = 8'h7e;
mem[7887] = 8'hd0;
mem[7888] = 8'hfe;
mem[7889] = 8'h68;
mem[7890] = 8'h48;
mem[7891] = 8'h09;
mem[7892] = 8'h08;
mem[7893] = 8'hc9;
mem[7894] = 8'hb8;
mem[7895] = 8'hd0;
mem[7896] = 8'hfe;
mem[7897] = 8'h28;
mem[7898] = 8'ha9;
mem[7899] = 8'hff;
mem[7900] = 8'h48;
mem[7901] = 8'ha2;
mem[7902] = 8'h80;
mem[7903] = 8'h28;
mem[7904] = 8'hec;
mem[7905] = 8'h1b;
mem[7906] = 8'h02;
mem[7907] = 8'h08;
mem[7908] = 8'h68;
mem[7909] = 8'h48;
mem[7910] = 8'h09;
mem[7911] = 8'h08;
mem[7912] = 8'hc9;
mem[7913] = 8'h7d;
mem[7914] = 8'hd0;
mem[7915] = 8'hfe;
mem[7916] = 8'h28;
mem[7917] = 8'hca;
mem[7918] = 8'hec;
mem[7919] = 8'h1b;
mem[7920] = 8'h02;
mem[7921] = 8'h08;
mem[7922] = 8'h68;
mem[7923] = 8'h48;
mem[7924] = 8'h09;
mem[7925] = 8'h08;
mem[7926] = 8'hc9;
mem[7927] = 8'h7f;
mem[7928] = 8'hd0;
mem[7929] = 8'hfe;
mem[7930] = 8'h28;
mem[7931] = 8'hca;
mem[7932] = 8'hec;
mem[7933] = 8'h1b;
mem[7934] = 8'h02;
mem[7935] = 8'h08;
mem[7936] = 8'he0;
mem[7937] = 8'h7e;
mem[7938] = 8'hd0;
mem[7939] = 8'hfe;
mem[7940] = 8'h68;
mem[7941] = 8'h48;
mem[7942] = 8'h09;
mem[7943] = 8'h08;
mem[7944] = 8'hc9;
mem[7945] = 8'hfc;
mem[7946] = 8'hd0;
mem[7947] = 8'hfe;
mem[7948] = 8'h28;
mem[7949] = 8'ha9;
mem[7950] = 8'h00;
mem[7951] = 8'h48;
mem[7952] = 8'ha2;
mem[7953] = 8'h80;
mem[7954] = 8'h28;
mem[7955] = 8'he0;
mem[7956] = 8'h7f;
mem[7957] = 8'h08;
mem[7958] = 8'h68;
mem[7959] = 8'h48;
mem[7960] = 8'h09;
mem[7961] = 8'h08;
mem[7962] = 8'hc9;
mem[7963] = 8'h39;
mem[7964] = 8'hd0;
mem[7965] = 8'hfe;
mem[7966] = 8'h28;
mem[7967] = 8'hca;
mem[7968] = 8'he0;
mem[7969] = 8'h7f;
mem[7970] = 8'h08;
mem[7971] = 8'h68;
mem[7972] = 8'h48;
mem[7973] = 8'h09;
mem[7974] = 8'h08;
mem[7975] = 8'hc9;
mem[7976] = 8'h3b;
mem[7977] = 8'hd0;
mem[7978] = 8'hfe;
mem[7979] = 8'h28;
mem[7980] = 8'hca;
mem[7981] = 8'he0;
mem[7982] = 8'h7f;
mem[7983] = 8'h08;
mem[7984] = 8'he0;
mem[7985] = 8'h7e;
mem[7986] = 8'hd0;
mem[7987] = 8'hfe;
mem[7988] = 8'h68;
mem[7989] = 8'h48;
mem[7990] = 8'h09;
mem[7991] = 8'h08;
mem[7992] = 8'hc9;
mem[7993] = 8'hb8;
mem[7994] = 8'hd0;
mem[7995] = 8'hfe;
mem[7996] = 8'h28;
mem[7997] = 8'ha9;
mem[7998] = 8'hff;
mem[7999] = 8'h48;
mem[8000] = 8'ha2;
mem[8001] = 8'h80;
mem[8002] = 8'h28;
mem[8003] = 8'he0;
mem[8004] = 8'h7f;
mem[8005] = 8'h08;
mem[8006] = 8'h68;
mem[8007] = 8'h48;
mem[8008] = 8'h09;
mem[8009] = 8'h08;
mem[8010] = 8'hc9;
mem[8011] = 8'h7d;
mem[8012] = 8'hd0;
mem[8013] = 8'hfe;
mem[8014] = 8'h28;
mem[8015] = 8'hca;
mem[8016] = 8'he0;
mem[8017] = 8'h7f;
mem[8018] = 8'h08;
mem[8019] = 8'h68;
mem[8020] = 8'h48;
mem[8021] = 8'h09;
mem[8022] = 8'h08;
mem[8023] = 8'hc9;
mem[8024] = 8'h7f;
mem[8025] = 8'hd0;
mem[8026] = 8'hfe;
mem[8027] = 8'h28;
mem[8028] = 8'hca;
mem[8029] = 8'he0;
mem[8030] = 8'h7f;
mem[8031] = 8'h08;
mem[8032] = 8'he0;
mem[8033] = 8'h7e;
mem[8034] = 8'hd0;
mem[8035] = 8'hfe;
mem[8036] = 8'h68;
mem[8037] = 8'h48;
mem[8038] = 8'h09;
mem[8039] = 8'h08;
mem[8040] = 8'hc9;
mem[8041] = 8'hfc;
mem[8042] = 8'hd0;
mem[8043] = 8'hfe;
mem[8044] = 8'h28;
mem[8045] = 8'had;
mem[8046] = 8'h00;
mem[8047] = 8'h02;
mem[8048] = 8'hc9;
mem[8049] = 8'h1a;
mem[8050] = 8'hd0;
mem[8051] = 8'hfe;
mem[8052] = 8'ha9;
mem[8053] = 8'h1b;
mem[8054] = 8'h8d;
mem[8055] = 8'h00;
mem[8056] = 8'h02;
mem[8057] = 8'ha9;
mem[8058] = 8'h00;
mem[8059] = 8'h48;
mem[8060] = 8'ha0;
mem[8061] = 8'h80;
mem[8062] = 8'h28;
mem[8063] = 8'hc4;
mem[8064] = 8'h17;
mem[8065] = 8'h08;
mem[8066] = 8'h68;
mem[8067] = 8'h48;
mem[8068] = 8'h09;
mem[8069] = 8'h08;
mem[8070] = 8'hc9;
mem[8071] = 8'h39;
mem[8072] = 8'hd0;
mem[8073] = 8'hfe;
mem[8074] = 8'h28;
mem[8075] = 8'h88;
mem[8076] = 8'hc4;
mem[8077] = 8'h17;
mem[8078] = 8'h08;
mem[8079] = 8'h68;
mem[8080] = 8'h48;
mem[8081] = 8'h09;
mem[8082] = 8'h08;
mem[8083] = 8'hc9;
mem[8084] = 8'h3b;
mem[8085] = 8'hd0;
mem[8086] = 8'hfe;
mem[8087] = 8'h28;
mem[8088] = 8'h88;
mem[8089] = 8'hc4;
mem[8090] = 8'h17;
mem[8091] = 8'h08;
mem[8092] = 8'hc0;
mem[8093] = 8'h7e;
mem[8094] = 8'hd0;
mem[8095] = 8'hfe;
mem[8096] = 8'h68;
mem[8097] = 8'h48;
mem[8098] = 8'h09;
mem[8099] = 8'h08;
mem[8100] = 8'hc9;
mem[8101] = 8'hb8;
mem[8102] = 8'hd0;
mem[8103] = 8'hfe;
mem[8104] = 8'h28;
mem[8105] = 8'ha9;
mem[8106] = 8'hff;
mem[8107] = 8'h48;
mem[8108] = 8'ha0;
mem[8109] = 8'h80;
mem[8110] = 8'h28;
mem[8111] = 8'hc4;
mem[8112] = 8'h17;
mem[8113] = 8'h08;
mem[8114] = 8'h68;
mem[8115] = 8'h48;
mem[8116] = 8'h09;
mem[8117] = 8'h08;
mem[8118] = 8'hc9;
mem[8119] = 8'h7d;
mem[8120] = 8'hd0;
mem[8121] = 8'hfe;
mem[8122] = 8'h28;
mem[8123] = 8'h88;
mem[8124] = 8'hc4;
mem[8125] = 8'h17;
mem[8126] = 8'h08;
mem[8127] = 8'h68;
mem[8128] = 8'h48;
mem[8129] = 8'h09;
mem[8130] = 8'h08;
mem[8131] = 8'hc9;
mem[8132] = 8'h7f;
mem[8133] = 8'hd0;
mem[8134] = 8'hfe;
mem[8135] = 8'h28;
mem[8136] = 8'h88;
mem[8137] = 8'hc4;
mem[8138] = 8'h17;
mem[8139] = 8'h08;
mem[8140] = 8'hc0;
mem[8141] = 8'h7e;
mem[8142] = 8'hd0;
mem[8143] = 8'hfe;
mem[8144] = 8'h68;
mem[8145] = 8'h48;
mem[8146] = 8'h09;
mem[8147] = 8'h08;
mem[8148] = 8'hc9;
mem[8149] = 8'hfc;
mem[8150] = 8'hd0;
mem[8151] = 8'hfe;
mem[8152] = 8'h28;
mem[8153] = 8'ha9;
mem[8154] = 8'h00;
mem[8155] = 8'h48;
mem[8156] = 8'ha0;
mem[8157] = 8'h80;
mem[8158] = 8'h28;
mem[8159] = 8'hcc;
mem[8160] = 8'h1b;
mem[8161] = 8'h02;
mem[8162] = 8'h08;
mem[8163] = 8'h68;
mem[8164] = 8'h48;
mem[8165] = 8'h09;
mem[8166] = 8'h08;
mem[8167] = 8'hc9;
mem[8168] = 8'h39;
mem[8169] = 8'hd0;
mem[8170] = 8'hfe;
mem[8171] = 8'h28;
mem[8172] = 8'h88;
mem[8173] = 8'hcc;
mem[8174] = 8'h1b;
mem[8175] = 8'h02;
mem[8176] = 8'h08;
mem[8177] = 8'h68;
mem[8178] = 8'h48;
mem[8179] = 8'h09;
mem[8180] = 8'h08;
mem[8181] = 8'hc9;
mem[8182] = 8'h3b;
mem[8183] = 8'hd0;
mem[8184] = 8'hfe;
mem[8185] = 8'h28;
mem[8186] = 8'h88;
mem[8187] = 8'hcc;
mem[8188] = 8'h1b;
mem[8189] = 8'h02;
mem[8190] = 8'h08;
mem[8191] = 8'hc0;
mem[8192] = 8'h7e;
mem[8193] = 8'hd0;
mem[8194] = 8'hfe;
mem[8195] = 8'h68;
mem[8196] = 8'h48;
mem[8197] = 8'h09;
mem[8198] = 8'h08;
mem[8199] = 8'hc9;
mem[8200] = 8'hb8;
mem[8201] = 8'hd0;
mem[8202] = 8'hfe;
mem[8203] = 8'h28;
mem[8204] = 8'ha9;
mem[8205] = 8'hff;
mem[8206] = 8'h48;
mem[8207] = 8'ha0;
mem[8208] = 8'h80;
mem[8209] = 8'h28;
mem[8210] = 8'hcc;
mem[8211] = 8'h1b;
mem[8212] = 8'h02;
mem[8213] = 8'h08;
mem[8214] = 8'h68;
mem[8215] = 8'h48;
mem[8216] = 8'h09;
mem[8217] = 8'h08;
mem[8218] = 8'hc9;
mem[8219] = 8'h7d;
mem[8220] = 8'hd0;
mem[8221] = 8'hfe;
mem[8222] = 8'h28;
mem[8223] = 8'h88;
mem[8224] = 8'hcc;
mem[8225] = 8'h1b;
mem[8226] = 8'h02;
mem[8227] = 8'h08;
mem[8228] = 8'h68;
mem[8229] = 8'h48;
mem[8230] = 8'h09;
mem[8231] = 8'h08;
mem[8232] = 8'hc9;
mem[8233] = 8'h7f;
mem[8234] = 8'hd0;
mem[8235] = 8'hfe;
mem[8236] = 8'h28;
mem[8237] = 8'h88;
mem[8238] = 8'hcc;
mem[8239] = 8'h1b;
mem[8240] = 8'h02;
mem[8241] = 8'h08;
mem[8242] = 8'hc0;
mem[8243] = 8'h7e;
mem[8244] = 8'hd0;
mem[8245] = 8'hfe;
mem[8246] = 8'h68;
mem[8247] = 8'h48;
mem[8248] = 8'h09;
mem[8249] = 8'h08;
mem[8250] = 8'hc9;
mem[8251] = 8'hfc;
mem[8252] = 8'hd0;
mem[8253] = 8'hfe;
mem[8254] = 8'h28;
mem[8255] = 8'ha9;
mem[8256] = 8'h00;
mem[8257] = 8'h48;
mem[8258] = 8'ha0;
mem[8259] = 8'h80;
mem[8260] = 8'h28;
mem[8261] = 8'hc0;
mem[8262] = 8'h7f;
mem[8263] = 8'h08;
mem[8264] = 8'h68;
mem[8265] = 8'h48;
mem[8266] = 8'h09;
mem[8267] = 8'h08;
mem[8268] = 8'hc9;
mem[8269] = 8'h39;
mem[8270] = 8'hd0;
mem[8271] = 8'hfe;
mem[8272] = 8'h28;
mem[8273] = 8'h88;
mem[8274] = 8'hc0;
mem[8275] = 8'h7f;
mem[8276] = 8'h08;
mem[8277] = 8'h68;
mem[8278] = 8'h48;
mem[8279] = 8'h09;
mem[8280] = 8'h08;
mem[8281] = 8'hc9;
mem[8282] = 8'h3b;
mem[8283] = 8'hd0;
mem[8284] = 8'hfe;
mem[8285] = 8'h28;
mem[8286] = 8'h88;
mem[8287] = 8'hc0;
mem[8288] = 8'h7f;
mem[8289] = 8'h08;
mem[8290] = 8'hc0;
mem[8291] = 8'h7e;
mem[8292] = 8'hd0;
mem[8293] = 8'hfe;
mem[8294] = 8'h68;
mem[8295] = 8'h48;
mem[8296] = 8'h09;
mem[8297] = 8'h08;
mem[8298] = 8'hc9;
mem[8299] = 8'hb8;
mem[8300] = 8'hd0;
mem[8301] = 8'hfe;
mem[8302] = 8'h28;
mem[8303] = 8'ha9;
mem[8304] = 8'hff;
mem[8305] = 8'h48;
mem[8306] = 8'ha0;
mem[8307] = 8'h80;
mem[8308] = 8'h28;
mem[8309] = 8'hc0;
mem[8310] = 8'h7f;
mem[8311] = 8'h08;
mem[8312] = 8'h68;
mem[8313] = 8'h48;
mem[8314] = 8'h09;
mem[8315] = 8'h08;
mem[8316] = 8'hc9;
mem[8317] = 8'h7d;
mem[8318] = 8'hd0;
mem[8319] = 8'hfe;
mem[8320] = 8'h28;
mem[8321] = 8'h88;
mem[8322] = 8'hc0;
mem[8323] = 8'h7f;
mem[8324] = 8'h08;
mem[8325] = 8'h68;
mem[8326] = 8'h48;
mem[8327] = 8'h09;
mem[8328] = 8'h08;
mem[8329] = 8'hc9;
mem[8330] = 8'h7f;
mem[8331] = 8'hd0;
mem[8332] = 8'hfe;
mem[8333] = 8'h28;
mem[8334] = 8'h88;
mem[8335] = 8'hc0;
mem[8336] = 8'h7f;
mem[8337] = 8'h08;
mem[8338] = 8'hc0;
mem[8339] = 8'h7e;
mem[8340] = 8'hd0;
mem[8341] = 8'hfe;
mem[8342] = 8'h68;
mem[8343] = 8'h48;
mem[8344] = 8'h09;
mem[8345] = 8'h08;
mem[8346] = 8'hc9;
mem[8347] = 8'hfc;
mem[8348] = 8'hd0;
mem[8349] = 8'hfe;
mem[8350] = 8'h28;
mem[8351] = 8'had;
mem[8352] = 8'h00;
mem[8353] = 8'h02;
mem[8354] = 8'hc9;
mem[8355] = 8'h1b;
mem[8356] = 8'hd0;
mem[8357] = 8'hfe;
mem[8358] = 8'ha9;
mem[8359] = 8'h1c;
mem[8360] = 8'h8d;
mem[8361] = 8'h00;
mem[8362] = 8'h02;
mem[8363] = 8'ha9;
mem[8364] = 8'h00;
mem[8365] = 8'h48;
mem[8366] = 8'ha9;
mem[8367] = 8'h80;
mem[8368] = 8'h28;
mem[8369] = 8'hc5;
mem[8370] = 8'h17;
mem[8371] = 8'h08;
mem[8372] = 8'hc9;
mem[8373] = 8'h80;
mem[8374] = 8'hd0;
mem[8375] = 8'hfe;
mem[8376] = 8'h68;
mem[8377] = 8'h48;
mem[8378] = 8'h09;
mem[8379] = 8'h08;
mem[8380] = 8'hc9;
mem[8381] = 8'h39;
mem[8382] = 8'hd0;
mem[8383] = 8'hfe;
mem[8384] = 8'h28;
mem[8385] = 8'ha9;
mem[8386] = 8'h00;
mem[8387] = 8'h48;
mem[8388] = 8'ha9;
mem[8389] = 8'h7f;
mem[8390] = 8'h28;
mem[8391] = 8'hc5;
mem[8392] = 8'h17;
mem[8393] = 8'h08;
mem[8394] = 8'hc9;
mem[8395] = 8'h7f;
mem[8396] = 8'hd0;
mem[8397] = 8'hfe;
mem[8398] = 8'h68;
mem[8399] = 8'h48;
mem[8400] = 8'h09;
mem[8401] = 8'h08;
mem[8402] = 8'hc9;
mem[8403] = 8'h3b;
mem[8404] = 8'hd0;
mem[8405] = 8'hfe;
mem[8406] = 8'h28;
mem[8407] = 8'ha9;
mem[8408] = 8'h00;
mem[8409] = 8'h48;
mem[8410] = 8'ha9;
mem[8411] = 8'h7e;
mem[8412] = 8'h28;
mem[8413] = 8'hc5;
mem[8414] = 8'h17;
mem[8415] = 8'h08;
mem[8416] = 8'hc9;
mem[8417] = 8'h7e;
mem[8418] = 8'hd0;
mem[8419] = 8'hfe;
mem[8420] = 8'h68;
mem[8421] = 8'h48;
mem[8422] = 8'h09;
mem[8423] = 8'h08;
mem[8424] = 8'hc9;
mem[8425] = 8'hb8;
mem[8426] = 8'hd0;
mem[8427] = 8'hfe;
mem[8428] = 8'h28;
mem[8429] = 8'ha9;
mem[8430] = 8'hff;
mem[8431] = 8'h48;
mem[8432] = 8'ha9;
mem[8433] = 8'h80;
mem[8434] = 8'h28;
mem[8435] = 8'hc5;
mem[8436] = 8'h17;
mem[8437] = 8'h08;
mem[8438] = 8'hc9;
mem[8439] = 8'h80;
mem[8440] = 8'hd0;
mem[8441] = 8'hfe;
mem[8442] = 8'h68;
mem[8443] = 8'h48;
mem[8444] = 8'h09;
mem[8445] = 8'h08;
mem[8446] = 8'hc9;
mem[8447] = 8'h7d;
mem[8448] = 8'hd0;
mem[8449] = 8'hfe;
mem[8450] = 8'h28;
mem[8451] = 8'ha9;
mem[8452] = 8'hff;
mem[8453] = 8'h48;
mem[8454] = 8'ha9;
mem[8455] = 8'h7f;
mem[8456] = 8'h28;
mem[8457] = 8'hc5;
mem[8458] = 8'h17;
mem[8459] = 8'h08;
mem[8460] = 8'hc9;
mem[8461] = 8'h7f;
mem[8462] = 8'hd0;
mem[8463] = 8'hfe;
mem[8464] = 8'h68;
mem[8465] = 8'h48;
mem[8466] = 8'h09;
mem[8467] = 8'h08;
mem[8468] = 8'hc9;
mem[8469] = 8'h7f;
mem[8470] = 8'hd0;
mem[8471] = 8'hfe;
mem[8472] = 8'h28;
mem[8473] = 8'ha9;
mem[8474] = 8'hff;
mem[8475] = 8'h48;
mem[8476] = 8'ha9;
mem[8477] = 8'h7e;
mem[8478] = 8'h28;
mem[8479] = 8'hc5;
mem[8480] = 8'h17;
mem[8481] = 8'h08;
mem[8482] = 8'hc9;
mem[8483] = 8'h7e;
mem[8484] = 8'hd0;
mem[8485] = 8'hfe;
mem[8486] = 8'h68;
mem[8487] = 8'h48;
mem[8488] = 8'h09;
mem[8489] = 8'h08;
mem[8490] = 8'hc9;
mem[8491] = 8'hfc;
mem[8492] = 8'hd0;
mem[8493] = 8'hfe;
mem[8494] = 8'h28;
mem[8495] = 8'ha9;
mem[8496] = 8'h00;
mem[8497] = 8'h48;
mem[8498] = 8'ha9;
mem[8499] = 8'h80;
mem[8500] = 8'h28;
mem[8501] = 8'hcd;
mem[8502] = 8'h1b;
mem[8503] = 8'h02;
mem[8504] = 8'h08;
mem[8505] = 8'hc9;
mem[8506] = 8'h80;
mem[8507] = 8'hd0;
mem[8508] = 8'hfe;
mem[8509] = 8'h68;
mem[8510] = 8'h48;
mem[8511] = 8'h09;
mem[8512] = 8'h08;
mem[8513] = 8'hc9;
mem[8514] = 8'h39;
mem[8515] = 8'hd0;
mem[8516] = 8'hfe;
mem[8517] = 8'h28;
mem[8518] = 8'ha9;
mem[8519] = 8'h00;
mem[8520] = 8'h48;
mem[8521] = 8'ha9;
mem[8522] = 8'h7f;
mem[8523] = 8'h28;
mem[8524] = 8'hcd;
mem[8525] = 8'h1b;
mem[8526] = 8'h02;
mem[8527] = 8'h08;
mem[8528] = 8'hc9;
mem[8529] = 8'h7f;
mem[8530] = 8'hd0;
mem[8531] = 8'hfe;
mem[8532] = 8'h68;
mem[8533] = 8'h48;
mem[8534] = 8'h09;
mem[8535] = 8'h08;
mem[8536] = 8'hc9;
mem[8537] = 8'h3b;
mem[8538] = 8'hd0;
mem[8539] = 8'hfe;
mem[8540] = 8'h28;
mem[8541] = 8'ha9;
mem[8542] = 8'h00;
mem[8543] = 8'h48;
mem[8544] = 8'ha9;
mem[8545] = 8'h7e;
mem[8546] = 8'h28;
mem[8547] = 8'hcd;
mem[8548] = 8'h1b;
mem[8549] = 8'h02;
mem[8550] = 8'h08;
mem[8551] = 8'hc9;
mem[8552] = 8'h7e;
mem[8553] = 8'hd0;
mem[8554] = 8'hfe;
mem[8555] = 8'h68;
mem[8556] = 8'h48;
mem[8557] = 8'h09;
mem[8558] = 8'h08;
mem[8559] = 8'hc9;
mem[8560] = 8'hb8;
mem[8561] = 8'hd0;
mem[8562] = 8'hfe;
mem[8563] = 8'h28;
mem[8564] = 8'ha9;
mem[8565] = 8'hff;
mem[8566] = 8'h48;
mem[8567] = 8'ha9;
mem[8568] = 8'h80;
mem[8569] = 8'h28;
mem[8570] = 8'hcd;
mem[8571] = 8'h1b;
mem[8572] = 8'h02;
mem[8573] = 8'h08;
mem[8574] = 8'hc9;
mem[8575] = 8'h80;
mem[8576] = 8'hd0;
mem[8577] = 8'hfe;
mem[8578] = 8'h68;
mem[8579] = 8'h48;
mem[8580] = 8'h09;
mem[8581] = 8'h08;
mem[8582] = 8'hc9;
mem[8583] = 8'h7d;
mem[8584] = 8'hd0;
mem[8585] = 8'hfe;
mem[8586] = 8'h28;
mem[8587] = 8'ha9;
mem[8588] = 8'hff;
mem[8589] = 8'h48;
mem[8590] = 8'ha9;
mem[8591] = 8'h7f;
mem[8592] = 8'h28;
mem[8593] = 8'hcd;
mem[8594] = 8'h1b;
mem[8595] = 8'h02;
mem[8596] = 8'h08;
mem[8597] = 8'hc9;
mem[8598] = 8'h7f;
mem[8599] = 8'hd0;
mem[8600] = 8'hfe;
mem[8601] = 8'h68;
mem[8602] = 8'h48;
mem[8603] = 8'h09;
mem[8604] = 8'h08;
mem[8605] = 8'hc9;
mem[8606] = 8'h7f;
mem[8607] = 8'hd0;
mem[8608] = 8'hfe;
mem[8609] = 8'h28;
mem[8610] = 8'ha9;
mem[8611] = 8'hff;
mem[8612] = 8'h48;
mem[8613] = 8'ha9;
mem[8614] = 8'h7e;
mem[8615] = 8'h28;
mem[8616] = 8'hcd;
mem[8617] = 8'h1b;
mem[8618] = 8'h02;
mem[8619] = 8'h08;
mem[8620] = 8'hc9;
mem[8621] = 8'h7e;
mem[8622] = 8'hd0;
mem[8623] = 8'hfe;
mem[8624] = 8'h68;
mem[8625] = 8'h48;
mem[8626] = 8'h09;
mem[8627] = 8'h08;
mem[8628] = 8'hc9;
mem[8629] = 8'hfc;
mem[8630] = 8'hd0;
mem[8631] = 8'hfe;
mem[8632] = 8'h28;
mem[8633] = 8'ha9;
mem[8634] = 8'h00;
mem[8635] = 8'h48;
mem[8636] = 8'ha9;
mem[8637] = 8'h80;
mem[8638] = 8'h28;
mem[8639] = 8'hc9;
mem[8640] = 8'h7f;
mem[8641] = 8'h08;
mem[8642] = 8'hc9;
mem[8643] = 8'h80;
mem[8644] = 8'hd0;
mem[8645] = 8'hfe;
mem[8646] = 8'h68;
mem[8647] = 8'h48;
mem[8648] = 8'h09;
mem[8649] = 8'h08;
mem[8650] = 8'hc9;
mem[8651] = 8'h39;
mem[8652] = 8'hd0;
mem[8653] = 8'hfe;
mem[8654] = 8'h28;
mem[8655] = 8'ha9;
mem[8656] = 8'h00;
mem[8657] = 8'h48;
mem[8658] = 8'ha9;
mem[8659] = 8'h7f;
mem[8660] = 8'h28;
mem[8661] = 8'hc9;
mem[8662] = 8'h7f;
mem[8663] = 8'h08;
mem[8664] = 8'hc9;
mem[8665] = 8'h7f;
mem[8666] = 8'hd0;
mem[8667] = 8'hfe;
mem[8668] = 8'h68;
mem[8669] = 8'h48;
mem[8670] = 8'h09;
mem[8671] = 8'h08;
mem[8672] = 8'hc9;
mem[8673] = 8'h3b;
mem[8674] = 8'hd0;
mem[8675] = 8'hfe;
mem[8676] = 8'h28;
mem[8677] = 8'ha9;
mem[8678] = 8'h00;
mem[8679] = 8'h48;
mem[8680] = 8'ha9;
mem[8681] = 8'h7e;
mem[8682] = 8'h28;
mem[8683] = 8'hc9;
mem[8684] = 8'h7f;
mem[8685] = 8'h08;
mem[8686] = 8'hc9;
mem[8687] = 8'h7e;
mem[8688] = 8'hd0;
mem[8689] = 8'hfe;
mem[8690] = 8'h68;
mem[8691] = 8'h48;
mem[8692] = 8'h09;
mem[8693] = 8'h08;
mem[8694] = 8'hc9;
mem[8695] = 8'hb8;
mem[8696] = 8'hd0;
mem[8697] = 8'hfe;
mem[8698] = 8'h28;
mem[8699] = 8'ha9;
mem[8700] = 8'hff;
mem[8701] = 8'h48;
mem[8702] = 8'ha9;
mem[8703] = 8'h80;
mem[8704] = 8'h28;
mem[8705] = 8'hc9;
mem[8706] = 8'h7f;
mem[8707] = 8'h08;
mem[8708] = 8'hc9;
mem[8709] = 8'h80;
mem[8710] = 8'hd0;
mem[8711] = 8'hfe;
mem[8712] = 8'h68;
mem[8713] = 8'h48;
mem[8714] = 8'h09;
mem[8715] = 8'h08;
mem[8716] = 8'hc9;
mem[8717] = 8'h7d;
mem[8718] = 8'hd0;
mem[8719] = 8'hfe;
mem[8720] = 8'h28;
mem[8721] = 8'ha9;
mem[8722] = 8'hff;
mem[8723] = 8'h48;
mem[8724] = 8'ha9;
mem[8725] = 8'h7f;
mem[8726] = 8'h28;
mem[8727] = 8'hc9;
mem[8728] = 8'h7f;
mem[8729] = 8'h08;
mem[8730] = 8'hc9;
mem[8731] = 8'h7f;
mem[8732] = 8'hd0;
mem[8733] = 8'hfe;
mem[8734] = 8'h68;
mem[8735] = 8'h48;
mem[8736] = 8'h09;
mem[8737] = 8'h08;
mem[8738] = 8'hc9;
mem[8739] = 8'h7f;
mem[8740] = 8'hd0;
mem[8741] = 8'hfe;
mem[8742] = 8'h28;
mem[8743] = 8'ha9;
mem[8744] = 8'hff;
mem[8745] = 8'h48;
mem[8746] = 8'ha9;
mem[8747] = 8'h7e;
mem[8748] = 8'h28;
mem[8749] = 8'hc9;
mem[8750] = 8'h7f;
mem[8751] = 8'h08;
mem[8752] = 8'hc9;
mem[8753] = 8'h7e;
mem[8754] = 8'hd0;
mem[8755] = 8'hfe;
mem[8756] = 8'h68;
mem[8757] = 8'h48;
mem[8758] = 8'h09;
mem[8759] = 8'h08;
mem[8760] = 8'hc9;
mem[8761] = 8'hfc;
mem[8762] = 8'hd0;
mem[8763] = 8'hfe;
mem[8764] = 8'h28;
mem[8765] = 8'ha2;
mem[8766] = 8'h04;
mem[8767] = 8'ha9;
mem[8768] = 8'h00;
mem[8769] = 8'h48;
mem[8770] = 8'ha9;
mem[8771] = 8'h80;
mem[8772] = 8'h28;
mem[8773] = 8'hd5;
mem[8774] = 8'h13;
mem[8775] = 8'h08;
mem[8776] = 8'hc9;
mem[8777] = 8'h80;
mem[8778] = 8'hd0;
mem[8779] = 8'hfe;
mem[8780] = 8'h68;
mem[8781] = 8'h48;
mem[8782] = 8'h09;
mem[8783] = 8'h08;
mem[8784] = 8'hc9;
mem[8785] = 8'h39;
mem[8786] = 8'hd0;
mem[8787] = 8'hfe;
mem[8788] = 8'h28;
mem[8789] = 8'ha9;
mem[8790] = 8'h00;
mem[8791] = 8'h48;
mem[8792] = 8'ha9;
mem[8793] = 8'h7f;
mem[8794] = 8'h28;
mem[8795] = 8'hd5;
mem[8796] = 8'h13;
mem[8797] = 8'h08;
mem[8798] = 8'hc9;
mem[8799] = 8'h7f;
mem[8800] = 8'hd0;
mem[8801] = 8'hfe;
mem[8802] = 8'h68;
mem[8803] = 8'h48;
mem[8804] = 8'h09;
mem[8805] = 8'h08;
mem[8806] = 8'hc9;
mem[8807] = 8'h3b;
mem[8808] = 8'hd0;
mem[8809] = 8'hfe;
mem[8810] = 8'h28;
mem[8811] = 8'ha9;
mem[8812] = 8'h00;
mem[8813] = 8'h48;
mem[8814] = 8'ha9;
mem[8815] = 8'h7e;
mem[8816] = 8'h28;
mem[8817] = 8'hd5;
mem[8818] = 8'h13;
mem[8819] = 8'h08;
mem[8820] = 8'hc9;
mem[8821] = 8'h7e;
mem[8822] = 8'hd0;
mem[8823] = 8'hfe;
mem[8824] = 8'h68;
mem[8825] = 8'h48;
mem[8826] = 8'h09;
mem[8827] = 8'h08;
mem[8828] = 8'hc9;
mem[8829] = 8'hb8;
mem[8830] = 8'hd0;
mem[8831] = 8'hfe;
mem[8832] = 8'h28;
mem[8833] = 8'ha9;
mem[8834] = 8'hff;
mem[8835] = 8'h48;
mem[8836] = 8'ha9;
mem[8837] = 8'h80;
mem[8838] = 8'h28;
mem[8839] = 8'hd5;
mem[8840] = 8'h13;
mem[8841] = 8'h08;
mem[8842] = 8'hc9;
mem[8843] = 8'h80;
mem[8844] = 8'hd0;
mem[8845] = 8'hfe;
mem[8846] = 8'h68;
mem[8847] = 8'h48;
mem[8848] = 8'h09;
mem[8849] = 8'h08;
mem[8850] = 8'hc9;
mem[8851] = 8'h7d;
mem[8852] = 8'hd0;
mem[8853] = 8'hfe;
mem[8854] = 8'h28;
mem[8855] = 8'ha9;
mem[8856] = 8'hff;
mem[8857] = 8'h48;
mem[8858] = 8'ha9;
mem[8859] = 8'h7f;
mem[8860] = 8'h28;
mem[8861] = 8'hd5;
mem[8862] = 8'h13;
mem[8863] = 8'h08;
mem[8864] = 8'hc9;
mem[8865] = 8'h7f;
mem[8866] = 8'hd0;
mem[8867] = 8'hfe;
mem[8868] = 8'h68;
mem[8869] = 8'h48;
mem[8870] = 8'h09;
mem[8871] = 8'h08;
mem[8872] = 8'hc9;
mem[8873] = 8'h7f;
mem[8874] = 8'hd0;
mem[8875] = 8'hfe;
mem[8876] = 8'h28;
mem[8877] = 8'ha9;
mem[8878] = 8'hff;
mem[8879] = 8'h48;
mem[8880] = 8'ha9;
mem[8881] = 8'h7e;
mem[8882] = 8'h28;
mem[8883] = 8'hd5;
mem[8884] = 8'h13;
mem[8885] = 8'h08;
mem[8886] = 8'hc9;
mem[8887] = 8'h7e;
mem[8888] = 8'hd0;
mem[8889] = 8'hfe;
mem[8890] = 8'h68;
mem[8891] = 8'h48;
mem[8892] = 8'h09;
mem[8893] = 8'h08;
mem[8894] = 8'hc9;
mem[8895] = 8'hfc;
mem[8896] = 8'hd0;
mem[8897] = 8'hfe;
mem[8898] = 8'h28;
mem[8899] = 8'ha9;
mem[8900] = 8'h00;
mem[8901] = 8'h48;
mem[8902] = 8'ha9;
mem[8903] = 8'h80;
mem[8904] = 8'h28;
mem[8905] = 8'hdd;
mem[8906] = 8'h17;
mem[8907] = 8'h02;
mem[8908] = 8'h08;
mem[8909] = 8'hc9;
mem[8910] = 8'h80;
mem[8911] = 8'hd0;
mem[8912] = 8'hfe;
mem[8913] = 8'h68;
mem[8914] = 8'h48;
mem[8915] = 8'h09;
mem[8916] = 8'h08;
mem[8917] = 8'hc9;
mem[8918] = 8'h39;
mem[8919] = 8'hd0;
mem[8920] = 8'hfe;
mem[8921] = 8'h28;
mem[8922] = 8'ha9;
mem[8923] = 8'h00;
mem[8924] = 8'h48;
mem[8925] = 8'ha9;
mem[8926] = 8'h7f;
mem[8927] = 8'h28;
mem[8928] = 8'hdd;
mem[8929] = 8'h17;
mem[8930] = 8'h02;
mem[8931] = 8'h08;
mem[8932] = 8'hc9;
mem[8933] = 8'h7f;
mem[8934] = 8'hd0;
mem[8935] = 8'hfe;
mem[8936] = 8'h68;
mem[8937] = 8'h48;
mem[8938] = 8'h09;
mem[8939] = 8'h08;
mem[8940] = 8'hc9;
mem[8941] = 8'h3b;
mem[8942] = 8'hd0;
mem[8943] = 8'hfe;
mem[8944] = 8'h28;
mem[8945] = 8'ha9;
mem[8946] = 8'h00;
mem[8947] = 8'h48;
mem[8948] = 8'ha9;
mem[8949] = 8'h7e;
mem[8950] = 8'h28;
mem[8951] = 8'hdd;
mem[8952] = 8'h17;
mem[8953] = 8'h02;
mem[8954] = 8'h08;
mem[8955] = 8'hc9;
mem[8956] = 8'h7e;
mem[8957] = 8'hd0;
mem[8958] = 8'hfe;
mem[8959] = 8'h68;
mem[8960] = 8'h48;
mem[8961] = 8'h09;
mem[8962] = 8'h08;
mem[8963] = 8'hc9;
mem[8964] = 8'hb8;
mem[8965] = 8'hd0;
mem[8966] = 8'hfe;
mem[8967] = 8'h28;
mem[8968] = 8'ha9;
mem[8969] = 8'hff;
mem[8970] = 8'h48;
mem[8971] = 8'ha9;
mem[8972] = 8'h80;
mem[8973] = 8'h28;
mem[8974] = 8'hdd;
mem[8975] = 8'h17;
mem[8976] = 8'h02;
mem[8977] = 8'h08;
mem[8978] = 8'hc9;
mem[8979] = 8'h80;
mem[8980] = 8'hd0;
mem[8981] = 8'hfe;
mem[8982] = 8'h68;
mem[8983] = 8'h48;
mem[8984] = 8'h09;
mem[8985] = 8'h08;
mem[8986] = 8'hc9;
mem[8987] = 8'h7d;
mem[8988] = 8'hd0;
mem[8989] = 8'hfe;
mem[8990] = 8'h28;
mem[8991] = 8'ha9;
mem[8992] = 8'hff;
mem[8993] = 8'h48;
mem[8994] = 8'ha9;
mem[8995] = 8'h7f;
mem[8996] = 8'h28;
mem[8997] = 8'hdd;
mem[8998] = 8'h17;
mem[8999] = 8'h02;
mem[9000] = 8'h08;
mem[9001] = 8'hc9;
mem[9002] = 8'h7f;
mem[9003] = 8'hd0;
mem[9004] = 8'hfe;
mem[9005] = 8'h68;
mem[9006] = 8'h48;
mem[9007] = 8'h09;
mem[9008] = 8'h08;
mem[9009] = 8'hc9;
mem[9010] = 8'h7f;
mem[9011] = 8'hd0;
mem[9012] = 8'hfe;
mem[9013] = 8'h28;
mem[9014] = 8'ha9;
mem[9015] = 8'hff;
mem[9016] = 8'h48;
mem[9017] = 8'ha9;
mem[9018] = 8'h7e;
mem[9019] = 8'h28;
mem[9020] = 8'hdd;
mem[9021] = 8'h17;
mem[9022] = 8'h02;
mem[9023] = 8'h08;
mem[9024] = 8'hc9;
mem[9025] = 8'h7e;
mem[9026] = 8'hd0;
mem[9027] = 8'hfe;
mem[9028] = 8'h68;
mem[9029] = 8'h48;
mem[9030] = 8'h09;
mem[9031] = 8'h08;
mem[9032] = 8'hc9;
mem[9033] = 8'hfc;
mem[9034] = 8'hd0;
mem[9035] = 8'hfe;
mem[9036] = 8'h28;
mem[9037] = 8'ha0;
mem[9038] = 8'h04;
mem[9039] = 8'ha2;
mem[9040] = 8'h08;
mem[9041] = 8'ha9;
mem[9042] = 8'h00;
mem[9043] = 8'h48;
mem[9044] = 8'ha9;
mem[9045] = 8'h80;
mem[9046] = 8'h28;
mem[9047] = 8'hd9;
mem[9048] = 8'h17;
mem[9049] = 8'h02;
mem[9050] = 8'h08;
mem[9051] = 8'hc9;
mem[9052] = 8'h80;
mem[9053] = 8'hd0;
mem[9054] = 8'hfe;
mem[9055] = 8'h68;
mem[9056] = 8'h48;
mem[9057] = 8'h09;
mem[9058] = 8'h08;
mem[9059] = 8'hc9;
mem[9060] = 8'h39;
mem[9061] = 8'hd0;
mem[9062] = 8'hfe;
mem[9063] = 8'h28;
mem[9064] = 8'ha9;
mem[9065] = 8'h00;
mem[9066] = 8'h48;
mem[9067] = 8'ha9;
mem[9068] = 8'h7f;
mem[9069] = 8'h28;
mem[9070] = 8'hd9;
mem[9071] = 8'h17;
mem[9072] = 8'h02;
mem[9073] = 8'h08;
mem[9074] = 8'hc9;
mem[9075] = 8'h7f;
mem[9076] = 8'hd0;
mem[9077] = 8'hfe;
mem[9078] = 8'h68;
mem[9079] = 8'h48;
mem[9080] = 8'h09;
mem[9081] = 8'h08;
mem[9082] = 8'hc9;
mem[9083] = 8'h3b;
mem[9084] = 8'hd0;
mem[9085] = 8'hfe;
mem[9086] = 8'h28;
mem[9087] = 8'ha9;
mem[9088] = 8'h00;
mem[9089] = 8'h48;
mem[9090] = 8'ha9;
mem[9091] = 8'h7e;
mem[9092] = 8'h28;
mem[9093] = 8'hd9;
mem[9094] = 8'h17;
mem[9095] = 8'h02;
mem[9096] = 8'h08;
mem[9097] = 8'hc9;
mem[9098] = 8'h7e;
mem[9099] = 8'hd0;
mem[9100] = 8'hfe;
mem[9101] = 8'h68;
mem[9102] = 8'h48;
mem[9103] = 8'h09;
mem[9104] = 8'h08;
mem[9105] = 8'hc9;
mem[9106] = 8'hb8;
mem[9107] = 8'hd0;
mem[9108] = 8'hfe;
mem[9109] = 8'h28;
mem[9110] = 8'ha9;
mem[9111] = 8'hff;
mem[9112] = 8'h48;
mem[9113] = 8'ha9;
mem[9114] = 8'h80;
mem[9115] = 8'h28;
mem[9116] = 8'hd9;
mem[9117] = 8'h17;
mem[9118] = 8'h02;
mem[9119] = 8'h08;
mem[9120] = 8'hc9;
mem[9121] = 8'h80;
mem[9122] = 8'hd0;
mem[9123] = 8'hfe;
mem[9124] = 8'h68;
mem[9125] = 8'h48;
mem[9126] = 8'h09;
mem[9127] = 8'h08;
mem[9128] = 8'hc9;
mem[9129] = 8'h7d;
mem[9130] = 8'hd0;
mem[9131] = 8'hfe;
mem[9132] = 8'h28;
mem[9133] = 8'ha9;
mem[9134] = 8'hff;
mem[9135] = 8'h48;
mem[9136] = 8'ha9;
mem[9137] = 8'h7f;
mem[9138] = 8'h28;
mem[9139] = 8'hd9;
mem[9140] = 8'h17;
mem[9141] = 8'h02;
mem[9142] = 8'h08;
mem[9143] = 8'hc9;
mem[9144] = 8'h7f;
mem[9145] = 8'hd0;
mem[9146] = 8'hfe;
mem[9147] = 8'h68;
mem[9148] = 8'h48;
mem[9149] = 8'h09;
mem[9150] = 8'h08;
mem[9151] = 8'hc9;
mem[9152] = 8'h7f;
mem[9153] = 8'hd0;
mem[9154] = 8'hfe;
mem[9155] = 8'h28;
mem[9156] = 8'ha9;
mem[9157] = 8'hff;
mem[9158] = 8'h48;
mem[9159] = 8'ha9;
mem[9160] = 8'h7e;
mem[9161] = 8'h28;
mem[9162] = 8'hd9;
mem[9163] = 8'h17;
mem[9164] = 8'h02;
mem[9165] = 8'h08;
mem[9166] = 8'hc9;
mem[9167] = 8'h7e;
mem[9168] = 8'hd0;
mem[9169] = 8'hfe;
mem[9170] = 8'h68;
mem[9171] = 8'h48;
mem[9172] = 8'h09;
mem[9173] = 8'h08;
mem[9174] = 8'hc9;
mem[9175] = 8'hfc;
mem[9176] = 8'hd0;
mem[9177] = 8'hfe;
mem[9178] = 8'h28;
mem[9179] = 8'ha9;
mem[9180] = 8'h00;
mem[9181] = 8'h48;
mem[9182] = 8'ha9;
mem[9183] = 8'h80;
mem[9184] = 8'h28;
mem[9185] = 8'hc1;
mem[9186] = 8'h24;
mem[9187] = 8'h08;
mem[9188] = 8'hc9;
mem[9189] = 8'h80;
mem[9190] = 8'hd0;
mem[9191] = 8'hfe;
mem[9192] = 8'h68;
mem[9193] = 8'h48;
mem[9194] = 8'h09;
mem[9195] = 8'h08;
mem[9196] = 8'hc9;
mem[9197] = 8'h39;
mem[9198] = 8'hd0;
mem[9199] = 8'hfe;
mem[9200] = 8'h28;
mem[9201] = 8'ha9;
mem[9202] = 8'h00;
mem[9203] = 8'h48;
mem[9204] = 8'ha9;
mem[9205] = 8'h7f;
mem[9206] = 8'h28;
mem[9207] = 8'hc1;
mem[9208] = 8'h24;
mem[9209] = 8'h08;
mem[9210] = 8'hc9;
mem[9211] = 8'h7f;
mem[9212] = 8'hd0;
mem[9213] = 8'hfe;
mem[9214] = 8'h68;
mem[9215] = 8'h48;
mem[9216] = 8'h09;
mem[9217] = 8'h08;
mem[9218] = 8'hc9;
mem[9219] = 8'h3b;
mem[9220] = 8'hd0;
mem[9221] = 8'hfe;
mem[9222] = 8'h28;
mem[9223] = 8'ha9;
mem[9224] = 8'h00;
mem[9225] = 8'h48;
mem[9226] = 8'ha9;
mem[9227] = 8'h7e;
mem[9228] = 8'h28;
mem[9229] = 8'hc1;
mem[9230] = 8'h24;
mem[9231] = 8'h08;
mem[9232] = 8'hc9;
mem[9233] = 8'h7e;
mem[9234] = 8'hd0;
mem[9235] = 8'hfe;
mem[9236] = 8'h68;
mem[9237] = 8'h48;
mem[9238] = 8'h09;
mem[9239] = 8'h08;
mem[9240] = 8'hc9;
mem[9241] = 8'hb8;
mem[9242] = 8'hd0;
mem[9243] = 8'hfe;
mem[9244] = 8'h28;
mem[9245] = 8'ha9;
mem[9246] = 8'hff;
mem[9247] = 8'h48;
mem[9248] = 8'ha9;
mem[9249] = 8'h80;
mem[9250] = 8'h28;
mem[9251] = 8'hc1;
mem[9252] = 8'h24;
mem[9253] = 8'h08;
mem[9254] = 8'hc9;
mem[9255] = 8'h80;
mem[9256] = 8'hd0;
mem[9257] = 8'hfe;
mem[9258] = 8'h68;
mem[9259] = 8'h48;
mem[9260] = 8'h09;
mem[9261] = 8'h08;
mem[9262] = 8'hc9;
mem[9263] = 8'h7d;
mem[9264] = 8'hd0;
mem[9265] = 8'hfe;
mem[9266] = 8'h28;
mem[9267] = 8'ha9;
mem[9268] = 8'hff;
mem[9269] = 8'h48;
mem[9270] = 8'ha9;
mem[9271] = 8'h7f;
mem[9272] = 8'h28;
mem[9273] = 8'hc1;
mem[9274] = 8'h24;
mem[9275] = 8'h08;
mem[9276] = 8'hc9;
mem[9277] = 8'h7f;
mem[9278] = 8'hd0;
mem[9279] = 8'hfe;
mem[9280] = 8'h68;
mem[9281] = 8'h48;
mem[9282] = 8'h09;
mem[9283] = 8'h08;
mem[9284] = 8'hc9;
mem[9285] = 8'h7f;
mem[9286] = 8'hd0;
mem[9287] = 8'hfe;
mem[9288] = 8'h28;
mem[9289] = 8'ha9;
mem[9290] = 8'hff;
mem[9291] = 8'h48;
mem[9292] = 8'ha9;
mem[9293] = 8'h7e;
mem[9294] = 8'h28;
mem[9295] = 8'hc1;
mem[9296] = 8'h24;
mem[9297] = 8'h08;
mem[9298] = 8'hc9;
mem[9299] = 8'h7e;
mem[9300] = 8'hd0;
mem[9301] = 8'hfe;
mem[9302] = 8'h68;
mem[9303] = 8'h48;
mem[9304] = 8'h09;
mem[9305] = 8'h08;
mem[9306] = 8'hc9;
mem[9307] = 8'hfc;
mem[9308] = 8'hd0;
mem[9309] = 8'hfe;
mem[9310] = 8'h28;
mem[9311] = 8'ha9;
mem[9312] = 8'h00;
mem[9313] = 8'h48;
mem[9314] = 8'ha9;
mem[9315] = 8'h80;
mem[9316] = 8'h28;
mem[9317] = 8'hd1;
mem[9318] = 8'h24;
mem[9319] = 8'h08;
mem[9320] = 8'hc9;
mem[9321] = 8'h80;
mem[9322] = 8'hd0;
mem[9323] = 8'hfe;
mem[9324] = 8'h68;
mem[9325] = 8'h48;
mem[9326] = 8'h09;
mem[9327] = 8'h08;
mem[9328] = 8'hc9;
mem[9329] = 8'h39;
mem[9330] = 8'hd0;
mem[9331] = 8'hfe;
mem[9332] = 8'h28;
mem[9333] = 8'ha9;
mem[9334] = 8'h00;
mem[9335] = 8'h48;
mem[9336] = 8'ha9;
mem[9337] = 8'h7f;
mem[9338] = 8'h28;
mem[9339] = 8'hd1;
mem[9340] = 8'h24;
mem[9341] = 8'h08;
mem[9342] = 8'hc9;
mem[9343] = 8'h7f;
mem[9344] = 8'hd0;
mem[9345] = 8'hfe;
mem[9346] = 8'h68;
mem[9347] = 8'h48;
mem[9348] = 8'h09;
mem[9349] = 8'h08;
mem[9350] = 8'hc9;
mem[9351] = 8'h3b;
mem[9352] = 8'hd0;
mem[9353] = 8'hfe;
mem[9354] = 8'h28;
mem[9355] = 8'ha9;
mem[9356] = 8'h00;
mem[9357] = 8'h48;
mem[9358] = 8'ha9;
mem[9359] = 8'h7e;
mem[9360] = 8'h28;
mem[9361] = 8'hd1;
mem[9362] = 8'h24;
mem[9363] = 8'h08;
mem[9364] = 8'hc9;
mem[9365] = 8'h7e;
mem[9366] = 8'hd0;
mem[9367] = 8'hfe;
mem[9368] = 8'h68;
mem[9369] = 8'h48;
mem[9370] = 8'h09;
mem[9371] = 8'h08;
mem[9372] = 8'hc9;
mem[9373] = 8'hb8;
mem[9374] = 8'hd0;
mem[9375] = 8'hfe;
mem[9376] = 8'h28;
mem[9377] = 8'ha9;
mem[9378] = 8'hff;
mem[9379] = 8'h48;
mem[9380] = 8'ha9;
mem[9381] = 8'h80;
mem[9382] = 8'h28;
mem[9383] = 8'hd1;
mem[9384] = 8'h24;
mem[9385] = 8'h08;
mem[9386] = 8'hc9;
mem[9387] = 8'h80;
mem[9388] = 8'hd0;
mem[9389] = 8'hfe;
mem[9390] = 8'h68;
mem[9391] = 8'h48;
mem[9392] = 8'h09;
mem[9393] = 8'h08;
mem[9394] = 8'hc9;
mem[9395] = 8'h7d;
mem[9396] = 8'hd0;
mem[9397] = 8'hfe;
mem[9398] = 8'h28;
mem[9399] = 8'ha9;
mem[9400] = 8'hff;
mem[9401] = 8'h48;
mem[9402] = 8'ha9;
mem[9403] = 8'h7f;
mem[9404] = 8'h28;
mem[9405] = 8'hd1;
mem[9406] = 8'h24;
mem[9407] = 8'h08;
mem[9408] = 8'hc9;
mem[9409] = 8'h7f;
mem[9410] = 8'hd0;
mem[9411] = 8'hfe;
mem[9412] = 8'h68;
mem[9413] = 8'h48;
mem[9414] = 8'h09;
mem[9415] = 8'h08;
mem[9416] = 8'hc9;
mem[9417] = 8'h7f;
mem[9418] = 8'hd0;
mem[9419] = 8'hfe;
mem[9420] = 8'h28;
mem[9421] = 8'ha9;
mem[9422] = 8'hff;
mem[9423] = 8'h48;
mem[9424] = 8'ha9;
mem[9425] = 8'h7e;
mem[9426] = 8'h28;
mem[9427] = 8'hd1;
mem[9428] = 8'h24;
mem[9429] = 8'h08;
mem[9430] = 8'hc9;
mem[9431] = 8'h7e;
mem[9432] = 8'hd0;
mem[9433] = 8'hfe;
mem[9434] = 8'h68;
mem[9435] = 8'h48;
mem[9436] = 8'h09;
mem[9437] = 8'h08;
mem[9438] = 8'hc9;
mem[9439] = 8'hfc;
mem[9440] = 8'hd0;
mem[9441] = 8'hfe;
mem[9442] = 8'h28;
mem[9443] = 8'had;
mem[9444] = 8'h00;
mem[9445] = 8'h02;
mem[9446] = 8'hc9;
mem[9447] = 8'h1c;
mem[9448] = 8'hd0;
mem[9449] = 8'hfe;
mem[9450] = 8'ha9;
mem[9451] = 8'h1d;
mem[9452] = 8'h8d;
mem[9453] = 8'h00;
mem[9454] = 8'h02;
mem[9455] = 8'ha2;
mem[9456] = 8'h03;
mem[9457] = 8'ha9;
mem[9458] = 8'h00;
mem[9459] = 8'h48;
mem[9460] = 8'hb5;
mem[9461] = 8'h13;
mem[9462] = 8'h28;
mem[9463] = 8'h0a;
mem[9464] = 8'h08;
mem[9465] = 8'hdd;
mem[9466] = 8'h20;
mem[9467] = 8'h02;
mem[9468] = 8'hd0;
mem[9469] = 8'hfe;
mem[9470] = 8'h68;
mem[9471] = 8'h09;
mem[9472] = 8'h08;
mem[9473] = 8'h49;
mem[9474] = 8'h38;
mem[9475] = 8'hdd;
mem[9476] = 8'h30;
mem[9477] = 8'h02;
mem[9478] = 8'hd0;
mem[9479] = 8'hfe;
mem[9480] = 8'hca;
mem[9481] = 8'h10;
mem[9482] = 8'he6;
mem[9483] = 8'ha2;
mem[9484] = 8'h03;
mem[9485] = 8'ha9;
mem[9486] = 8'hff;
mem[9487] = 8'h48;
mem[9488] = 8'hb5;
mem[9489] = 8'h13;
mem[9490] = 8'h28;
mem[9491] = 8'h0a;
mem[9492] = 8'h08;
mem[9493] = 8'hdd;
mem[9494] = 8'h20;
mem[9495] = 8'h02;
mem[9496] = 8'hd0;
mem[9497] = 8'hfe;
mem[9498] = 8'h68;
mem[9499] = 8'h09;
mem[9500] = 8'h08;
mem[9501] = 8'h49;
mem[9502] = 8'h7c;
mem[9503] = 8'hdd;
mem[9504] = 8'h30;
mem[9505] = 8'h02;
mem[9506] = 8'hd0;
mem[9507] = 8'hfe;
mem[9508] = 8'hca;
mem[9509] = 8'h10;
mem[9510] = 8'he6;
mem[9511] = 8'ha2;
mem[9512] = 8'h03;
mem[9513] = 8'ha9;
mem[9514] = 8'h00;
mem[9515] = 8'h48;
mem[9516] = 8'hb5;
mem[9517] = 8'h13;
mem[9518] = 8'h28;
mem[9519] = 8'h4a;
mem[9520] = 8'h08;
mem[9521] = 8'hdd;
mem[9522] = 8'h28;
mem[9523] = 8'h02;
mem[9524] = 8'hd0;
mem[9525] = 8'hfe;
mem[9526] = 8'h68;
mem[9527] = 8'h09;
mem[9528] = 8'h08;
mem[9529] = 8'h49;
mem[9530] = 8'h38;
mem[9531] = 8'hdd;
mem[9532] = 8'h38;
mem[9533] = 8'h02;
mem[9534] = 8'hd0;
mem[9535] = 8'hfe;
mem[9536] = 8'hca;
mem[9537] = 8'h10;
mem[9538] = 8'he6;
mem[9539] = 8'ha2;
mem[9540] = 8'h03;
mem[9541] = 8'ha9;
mem[9542] = 8'hff;
mem[9543] = 8'h48;
mem[9544] = 8'hb5;
mem[9545] = 8'h13;
mem[9546] = 8'h28;
mem[9547] = 8'h4a;
mem[9548] = 8'h08;
mem[9549] = 8'hdd;
mem[9550] = 8'h28;
mem[9551] = 8'h02;
mem[9552] = 8'hd0;
mem[9553] = 8'hfe;
mem[9554] = 8'h68;
mem[9555] = 8'h09;
mem[9556] = 8'h08;
mem[9557] = 8'h49;
mem[9558] = 8'h7c;
mem[9559] = 8'hdd;
mem[9560] = 8'h38;
mem[9561] = 8'h02;
mem[9562] = 8'hd0;
mem[9563] = 8'hfe;
mem[9564] = 8'hca;
mem[9565] = 8'h10;
mem[9566] = 8'he6;
mem[9567] = 8'ha2;
mem[9568] = 8'h03;
mem[9569] = 8'ha9;
mem[9570] = 8'h00;
mem[9571] = 8'h48;
mem[9572] = 8'hb5;
mem[9573] = 8'h13;
mem[9574] = 8'h28;
mem[9575] = 8'h2a;
mem[9576] = 8'h08;
mem[9577] = 8'hdd;
mem[9578] = 8'h20;
mem[9579] = 8'h02;
mem[9580] = 8'hd0;
mem[9581] = 8'hfe;
mem[9582] = 8'h68;
mem[9583] = 8'h09;
mem[9584] = 8'h08;
mem[9585] = 8'h49;
mem[9586] = 8'h38;
mem[9587] = 8'hdd;
mem[9588] = 8'h30;
mem[9589] = 8'h02;
mem[9590] = 8'hd0;
mem[9591] = 8'hfe;
mem[9592] = 8'hca;
mem[9593] = 8'h10;
mem[9594] = 8'he6;
mem[9595] = 8'ha2;
mem[9596] = 8'h03;
mem[9597] = 8'ha9;
mem[9598] = 8'hfe;
mem[9599] = 8'h48;
mem[9600] = 8'hb5;
mem[9601] = 8'h13;
mem[9602] = 8'h28;
mem[9603] = 8'h2a;
mem[9604] = 8'h08;
mem[9605] = 8'hdd;
mem[9606] = 8'h20;
mem[9607] = 8'h02;
mem[9608] = 8'hd0;
mem[9609] = 8'hfe;
mem[9610] = 8'h68;
mem[9611] = 8'h09;
mem[9612] = 8'h08;
mem[9613] = 8'h49;
mem[9614] = 8'h7c;
mem[9615] = 8'hdd;
mem[9616] = 8'h30;
mem[9617] = 8'h02;
mem[9618] = 8'hd0;
mem[9619] = 8'hfe;
mem[9620] = 8'hca;
mem[9621] = 8'h10;
mem[9622] = 8'he6;
mem[9623] = 8'ha2;
mem[9624] = 8'h03;
mem[9625] = 8'ha9;
mem[9626] = 8'h01;
mem[9627] = 8'h48;
mem[9628] = 8'hb5;
mem[9629] = 8'h13;
mem[9630] = 8'h28;
mem[9631] = 8'h2a;
mem[9632] = 8'h08;
mem[9633] = 8'hdd;
mem[9634] = 8'h24;
mem[9635] = 8'h02;
mem[9636] = 8'hd0;
mem[9637] = 8'hfe;
mem[9638] = 8'h68;
mem[9639] = 8'h09;
mem[9640] = 8'h08;
mem[9641] = 8'h49;
mem[9642] = 8'h38;
mem[9643] = 8'hdd;
mem[9644] = 8'h34;
mem[9645] = 8'h02;
mem[9646] = 8'hd0;
mem[9647] = 8'hfe;
mem[9648] = 8'hca;
mem[9649] = 8'h10;
mem[9650] = 8'he6;
mem[9651] = 8'ha2;
mem[9652] = 8'h03;
mem[9653] = 8'ha9;
mem[9654] = 8'hff;
mem[9655] = 8'h48;
mem[9656] = 8'hb5;
mem[9657] = 8'h13;
mem[9658] = 8'h28;
mem[9659] = 8'h2a;
mem[9660] = 8'h08;
mem[9661] = 8'hdd;
mem[9662] = 8'h24;
mem[9663] = 8'h02;
mem[9664] = 8'hd0;
mem[9665] = 8'hfe;
mem[9666] = 8'h68;
mem[9667] = 8'h09;
mem[9668] = 8'h08;
mem[9669] = 8'h49;
mem[9670] = 8'h7c;
mem[9671] = 8'hdd;
mem[9672] = 8'h34;
mem[9673] = 8'h02;
mem[9674] = 8'hd0;
mem[9675] = 8'hfe;
mem[9676] = 8'hca;
mem[9677] = 8'h10;
mem[9678] = 8'he6;
mem[9679] = 8'ha2;
mem[9680] = 8'h03;
mem[9681] = 8'ha9;
mem[9682] = 8'h00;
mem[9683] = 8'h48;
mem[9684] = 8'hb5;
mem[9685] = 8'h13;
mem[9686] = 8'h28;
mem[9687] = 8'h6a;
mem[9688] = 8'h08;
mem[9689] = 8'hdd;
mem[9690] = 8'h28;
mem[9691] = 8'h02;
mem[9692] = 8'hd0;
mem[9693] = 8'hfe;
mem[9694] = 8'h68;
mem[9695] = 8'h09;
mem[9696] = 8'h08;
mem[9697] = 8'h49;
mem[9698] = 8'h38;
mem[9699] = 8'hdd;
mem[9700] = 8'h38;
mem[9701] = 8'h02;
mem[9702] = 8'hd0;
mem[9703] = 8'hfe;
mem[9704] = 8'hca;
mem[9705] = 8'h10;
mem[9706] = 8'he6;
mem[9707] = 8'ha2;
mem[9708] = 8'h03;
mem[9709] = 8'ha9;
mem[9710] = 8'hfe;
mem[9711] = 8'h48;
mem[9712] = 8'hb5;
mem[9713] = 8'h13;
mem[9714] = 8'h28;
mem[9715] = 8'h6a;
mem[9716] = 8'h08;
mem[9717] = 8'hdd;
mem[9718] = 8'h28;
mem[9719] = 8'h02;
mem[9720] = 8'hd0;
mem[9721] = 8'hfe;
mem[9722] = 8'h68;
mem[9723] = 8'h09;
mem[9724] = 8'h08;
mem[9725] = 8'h49;
mem[9726] = 8'h7c;
mem[9727] = 8'hdd;
mem[9728] = 8'h38;
mem[9729] = 8'h02;
mem[9730] = 8'hd0;
mem[9731] = 8'hfe;
mem[9732] = 8'hca;
mem[9733] = 8'h10;
mem[9734] = 8'he6;
mem[9735] = 8'ha2;
mem[9736] = 8'h03;
mem[9737] = 8'ha9;
mem[9738] = 8'h01;
mem[9739] = 8'h48;
mem[9740] = 8'hb5;
mem[9741] = 8'h13;
mem[9742] = 8'h28;
mem[9743] = 8'h6a;
mem[9744] = 8'h08;
mem[9745] = 8'hdd;
mem[9746] = 8'h2c;
mem[9747] = 8'h02;
mem[9748] = 8'hd0;
mem[9749] = 8'hfe;
mem[9750] = 8'h68;
mem[9751] = 8'h09;
mem[9752] = 8'h08;
mem[9753] = 8'h49;
mem[9754] = 8'h38;
mem[9755] = 8'hdd;
mem[9756] = 8'h3c;
mem[9757] = 8'h02;
mem[9758] = 8'hd0;
mem[9759] = 8'hfe;
mem[9760] = 8'hca;
mem[9761] = 8'h10;
mem[9762] = 8'he6;
mem[9763] = 8'ha2;
mem[9764] = 8'h03;
mem[9765] = 8'ha9;
mem[9766] = 8'hff;
mem[9767] = 8'h48;
mem[9768] = 8'hb5;
mem[9769] = 8'h13;
mem[9770] = 8'h28;
mem[9771] = 8'h6a;
mem[9772] = 8'h08;
mem[9773] = 8'hdd;
mem[9774] = 8'h2c;
mem[9775] = 8'h02;
mem[9776] = 8'hd0;
mem[9777] = 8'hfe;
mem[9778] = 8'h68;
mem[9779] = 8'h09;
mem[9780] = 8'h08;
mem[9781] = 8'h49;
mem[9782] = 8'h7c;
mem[9783] = 8'hdd;
mem[9784] = 8'h3c;
mem[9785] = 8'h02;
mem[9786] = 8'hd0;
mem[9787] = 8'hfe;
mem[9788] = 8'hca;
mem[9789] = 8'h10;
mem[9790] = 8'he6;
mem[9791] = 8'had;
mem[9792] = 8'h00;
mem[9793] = 8'h02;
mem[9794] = 8'hc9;
mem[9795] = 8'h1d;
mem[9796] = 8'hd0;
mem[9797] = 8'hfe;
mem[9798] = 8'ha9;
mem[9799] = 8'h1e;
mem[9800] = 8'h8d;
mem[9801] = 8'h00;
mem[9802] = 8'h02;
mem[9803] = 8'ha2;
mem[9804] = 8'h03;
mem[9805] = 8'ha9;
mem[9806] = 8'h00;
mem[9807] = 8'h48;
mem[9808] = 8'hb5;
mem[9809] = 8'h13;
mem[9810] = 8'h85;
mem[9811] = 8'h0c;
mem[9812] = 8'h28;
mem[9813] = 8'h06;
mem[9814] = 8'h0c;
mem[9815] = 8'h08;
mem[9816] = 8'ha5;
mem[9817] = 8'h0c;
mem[9818] = 8'hdd;
mem[9819] = 8'h20;
mem[9820] = 8'h02;
mem[9821] = 8'hd0;
mem[9822] = 8'hfe;
mem[9823] = 8'h68;
mem[9824] = 8'h09;
mem[9825] = 8'h08;
mem[9826] = 8'h49;
mem[9827] = 8'h38;
mem[9828] = 8'hdd;
mem[9829] = 8'h30;
mem[9830] = 8'h02;
mem[9831] = 8'hd0;
mem[9832] = 8'hfe;
mem[9833] = 8'hca;
mem[9834] = 8'h10;
mem[9835] = 8'he1;
mem[9836] = 8'ha2;
mem[9837] = 8'h03;
mem[9838] = 8'ha9;
mem[9839] = 8'hff;
mem[9840] = 8'h48;
mem[9841] = 8'hb5;
mem[9842] = 8'h13;
mem[9843] = 8'h85;
mem[9844] = 8'h0c;
mem[9845] = 8'h28;
mem[9846] = 8'h06;
mem[9847] = 8'h0c;
mem[9848] = 8'h08;
mem[9849] = 8'ha5;
mem[9850] = 8'h0c;
mem[9851] = 8'hdd;
mem[9852] = 8'h20;
mem[9853] = 8'h02;
mem[9854] = 8'hd0;
mem[9855] = 8'hfe;
mem[9856] = 8'h68;
mem[9857] = 8'h09;
mem[9858] = 8'h08;
mem[9859] = 8'h49;
mem[9860] = 8'h7c;
mem[9861] = 8'hdd;
mem[9862] = 8'h30;
mem[9863] = 8'h02;
mem[9864] = 8'hd0;
mem[9865] = 8'hfe;
mem[9866] = 8'hca;
mem[9867] = 8'h10;
mem[9868] = 8'he1;
mem[9869] = 8'ha2;
mem[9870] = 8'h03;
mem[9871] = 8'ha9;
mem[9872] = 8'h00;
mem[9873] = 8'h48;
mem[9874] = 8'hb5;
mem[9875] = 8'h13;
mem[9876] = 8'h85;
mem[9877] = 8'h0c;
mem[9878] = 8'h28;
mem[9879] = 8'h46;
mem[9880] = 8'h0c;
mem[9881] = 8'h08;
mem[9882] = 8'ha5;
mem[9883] = 8'h0c;
mem[9884] = 8'hdd;
mem[9885] = 8'h28;
mem[9886] = 8'h02;
mem[9887] = 8'hd0;
mem[9888] = 8'hfe;
mem[9889] = 8'h68;
mem[9890] = 8'h09;
mem[9891] = 8'h08;
mem[9892] = 8'h49;
mem[9893] = 8'h38;
mem[9894] = 8'hdd;
mem[9895] = 8'h38;
mem[9896] = 8'h02;
mem[9897] = 8'hd0;
mem[9898] = 8'hfe;
mem[9899] = 8'hca;
mem[9900] = 8'h10;
mem[9901] = 8'he1;
mem[9902] = 8'ha2;
mem[9903] = 8'h03;
mem[9904] = 8'ha9;
mem[9905] = 8'hff;
mem[9906] = 8'h48;
mem[9907] = 8'hb5;
mem[9908] = 8'h13;
mem[9909] = 8'h85;
mem[9910] = 8'h0c;
mem[9911] = 8'h28;
mem[9912] = 8'h46;
mem[9913] = 8'h0c;
mem[9914] = 8'h08;
mem[9915] = 8'ha5;
mem[9916] = 8'h0c;
mem[9917] = 8'hdd;
mem[9918] = 8'h28;
mem[9919] = 8'h02;
mem[9920] = 8'hd0;
mem[9921] = 8'hfe;
mem[9922] = 8'h68;
mem[9923] = 8'h09;
mem[9924] = 8'h08;
mem[9925] = 8'h49;
mem[9926] = 8'h7c;
mem[9927] = 8'hdd;
mem[9928] = 8'h38;
mem[9929] = 8'h02;
mem[9930] = 8'hd0;
mem[9931] = 8'hfe;
mem[9932] = 8'hca;
mem[9933] = 8'h10;
mem[9934] = 8'he1;
mem[9935] = 8'ha2;
mem[9936] = 8'h03;
mem[9937] = 8'ha9;
mem[9938] = 8'h00;
mem[9939] = 8'h48;
mem[9940] = 8'hb5;
mem[9941] = 8'h13;
mem[9942] = 8'h85;
mem[9943] = 8'h0c;
mem[9944] = 8'h28;
mem[9945] = 8'h26;
mem[9946] = 8'h0c;
mem[9947] = 8'h08;
mem[9948] = 8'ha5;
mem[9949] = 8'h0c;
mem[9950] = 8'hdd;
mem[9951] = 8'h20;
mem[9952] = 8'h02;
mem[9953] = 8'hd0;
mem[9954] = 8'hfe;
mem[9955] = 8'h68;
mem[9956] = 8'h09;
mem[9957] = 8'h08;
mem[9958] = 8'h49;
mem[9959] = 8'h38;
mem[9960] = 8'hdd;
mem[9961] = 8'h30;
mem[9962] = 8'h02;
mem[9963] = 8'hd0;
mem[9964] = 8'hfe;
mem[9965] = 8'hca;
mem[9966] = 8'h10;
mem[9967] = 8'he1;
mem[9968] = 8'ha2;
mem[9969] = 8'h03;
mem[9970] = 8'ha9;
mem[9971] = 8'hfe;
mem[9972] = 8'h48;
mem[9973] = 8'hb5;
mem[9974] = 8'h13;
mem[9975] = 8'h85;
mem[9976] = 8'h0c;
mem[9977] = 8'h28;
mem[9978] = 8'h26;
mem[9979] = 8'h0c;
mem[9980] = 8'h08;
mem[9981] = 8'ha5;
mem[9982] = 8'h0c;
mem[9983] = 8'hdd;
mem[9984] = 8'h20;
mem[9985] = 8'h02;
mem[9986] = 8'hd0;
mem[9987] = 8'hfe;
mem[9988] = 8'h68;
mem[9989] = 8'h09;
mem[9990] = 8'h08;
mem[9991] = 8'h49;
mem[9992] = 8'h7c;
mem[9993] = 8'hdd;
mem[9994] = 8'h30;
mem[9995] = 8'h02;
mem[9996] = 8'hd0;
mem[9997] = 8'hfe;
mem[9998] = 8'hca;
mem[9999] = 8'h10;
mem[10000] = 8'he1;
mem[10001] = 8'ha2;
mem[10002] = 8'h03;
mem[10003] = 8'ha9;
mem[10004] = 8'h01;
mem[10005] = 8'h48;
mem[10006] = 8'hb5;
mem[10007] = 8'h13;
mem[10008] = 8'h85;
mem[10009] = 8'h0c;
mem[10010] = 8'h28;
mem[10011] = 8'h26;
mem[10012] = 8'h0c;
mem[10013] = 8'h08;
mem[10014] = 8'ha5;
mem[10015] = 8'h0c;
mem[10016] = 8'hdd;
mem[10017] = 8'h24;
mem[10018] = 8'h02;
mem[10019] = 8'hd0;
mem[10020] = 8'hfe;
mem[10021] = 8'h68;
mem[10022] = 8'h09;
mem[10023] = 8'h08;
mem[10024] = 8'h49;
mem[10025] = 8'h38;
mem[10026] = 8'hdd;
mem[10027] = 8'h34;
mem[10028] = 8'h02;
mem[10029] = 8'hd0;
mem[10030] = 8'hfe;
mem[10031] = 8'hca;
mem[10032] = 8'h10;
mem[10033] = 8'he1;
mem[10034] = 8'ha2;
mem[10035] = 8'h03;
mem[10036] = 8'ha9;
mem[10037] = 8'hff;
mem[10038] = 8'h48;
mem[10039] = 8'hb5;
mem[10040] = 8'h13;
mem[10041] = 8'h85;
mem[10042] = 8'h0c;
mem[10043] = 8'h28;
mem[10044] = 8'h26;
mem[10045] = 8'h0c;
mem[10046] = 8'h08;
mem[10047] = 8'ha5;
mem[10048] = 8'h0c;
mem[10049] = 8'hdd;
mem[10050] = 8'h24;
mem[10051] = 8'h02;
mem[10052] = 8'hd0;
mem[10053] = 8'hfe;
mem[10054] = 8'h68;
mem[10055] = 8'h09;
mem[10056] = 8'h08;
mem[10057] = 8'h49;
mem[10058] = 8'h7c;
mem[10059] = 8'hdd;
mem[10060] = 8'h34;
mem[10061] = 8'h02;
mem[10062] = 8'hd0;
mem[10063] = 8'hfe;
mem[10064] = 8'hca;
mem[10065] = 8'h10;
mem[10066] = 8'he1;
mem[10067] = 8'ha2;
mem[10068] = 8'h03;
mem[10069] = 8'ha9;
mem[10070] = 8'h00;
mem[10071] = 8'h48;
mem[10072] = 8'hb5;
mem[10073] = 8'h13;
mem[10074] = 8'h85;
mem[10075] = 8'h0c;
mem[10076] = 8'h28;
mem[10077] = 8'h66;
mem[10078] = 8'h0c;
mem[10079] = 8'h08;
mem[10080] = 8'ha5;
mem[10081] = 8'h0c;
mem[10082] = 8'hdd;
mem[10083] = 8'h28;
mem[10084] = 8'h02;
mem[10085] = 8'hd0;
mem[10086] = 8'hfe;
mem[10087] = 8'h68;
mem[10088] = 8'h09;
mem[10089] = 8'h08;
mem[10090] = 8'h49;
mem[10091] = 8'h38;
mem[10092] = 8'hdd;
mem[10093] = 8'h38;
mem[10094] = 8'h02;
mem[10095] = 8'hd0;
mem[10096] = 8'hfe;
mem[10097] = 8'hca;
mem[10098] = 8'h10;
mem[10099] = 8'he1;
mem[10100] = 8'ha2;
mem[10101] = 8'h03;
mem[10102] = 8'ha9;
mem[10103] = 8'hfe;
mem[10104] = 8'h48;
mem[10105] = 8'hb5;
mem[10106] = 8'h13;
mem[10107] = 8'h85;
mem[10108] = 8'h0c;
mem[10109] = 8'h28;
mem[10110] = 8'h66;
mem[10111] = 8'h0c;
mem[10112] = 8'h08;
mem[10113] = 8'ha5;
mem[10114] = 8'h0c;
mem[10115] = 8'hdd;
mem[10116] = 8'h28;
mem[10117] = 8'h02;
mem[10118] = 8'hd0;
mem[10119] = 8'hfe;
mem[10120] = 8'h68;
mem[10121] = 8'h09;
mem[10122] = 8'h08;
mem[10123] = 8'h49;
mem[10124] = 8'h7c;
mem[10125] = 8'hdd;
mem[10126] = 8'h38;
mem[10127] = 8'h02;
mem[10128] = 8'hd0;
mem[10129] = 8'hfe;
mem[10130] = 8'hca;
mem[10131] = 8'h10;
mem[10132] = 8'he1;
mem[10133] = 8'ha2;
mem[10134] = 8'h03;
mem[10135] = 8'ha9;
mem[10136] = 8'h01;
mem[10137] = 8'h48;
mem[10138] = 8'hb5;
mem[10139] = 8'h13;
mem[10140] = 8'h85;
mem[10141] = 8'h0c;
mem[10142] = 8'h28;
mem[10143] = 8'h66;
mem[10144] = 8'h0c;
mem[10145] = 8'h08;
mem[10146] = 8'ha5;
mem[10147] = 8'h0c;
mem[10148] = 8'hdd;
mem[10149] = 8'h2c;
mem[10150] = 8'h02;
mem[10151] = 8'hd0;
mem[10152] = 8'hfe;
mem[10153] = 8'h68;
mem[10154] = 8'h09;
mem[10155] = 8'h08;
mem[10156] = 8'h49;
mem[10157] = 8'h38;
mem[10158] = 8'hdd;
mem[10159] = 8'h3c;
mem[10160] = 8'h02;
mem[10161] = 8'hd0;
mem[10162] = 8'hfe;
mem[10163] = 8'hca;
mem[10164] = 8'h10;
mem[10165] = 8'he1;
mem[10166] = 8'ha2;
mem[10167] = 8'h03;
mem[10168] = 8'ha9;
mem[10169] = 8'hff;
mem[10170] = 8'h48;
mem[10171] = 8'hb5;
mem[10172] = 8'h13;
mem[10173] = 8'h85;
mem[10174] = 8'h0c;
mem[10175] = 8'h28;
mem[10176] = 8'h66;
mem[10177] = 8'h0c;
mem[10178] = 8'h08;
mem[10179] = 8'ha5;
mem[10180] = 8'h0c;
mem[10181] = 8'hdd;
mem[10182] = 8'h2c;
mem[10183] = 8'h02;
mem[10184] = 8'hd0;
mem[10185] = 8'hfe;
mem[10186] = 8'h68;
mem[10187] = 8'h09;
mem[10188] = 8'h08;
mem[10189] = 8'h49;
mem[10190] = 8'h7c;
mem[10191] = 8'hdd;
mem[10192] = 8'h3c;
mem[10193] = 8'h02;
mem[10194] = 8'hd0;
mem[10195] = 8'hfe;
mem[10196] = 8'hca;
mem[10197] = 8'h10;
mem[10198] = 8'he1;
mem[10199] = 8'had;
mem[10200] = 8'h00;
mem[10201] = 8'h02;
mem[10202] = 8'hc9;
mem[10203] = 8'h1e;
mem[10204] = 8'hd0;
mem[10205] = 8'hfe;
mem[10206] = 8'ha9;
mem[10207] = 8'h1f;
mem[10208] = 8'h8d;
mem[10209] = 8'h00;
mem[10210] = 8'h02;
mem[10211] = 8'ha2;
mem[10212] = 8'h03;
mem[10213] = 8'ha9;
mem[10214] = 8'h00;
mem[10215] = 8'h48;
mem[10216] = 8'hb5;
mem[10217] = 8'h13;
mem[10218] = 8'h8d;
mem[10219] = 8'h03;
mem[10220] = 8'h02;
mem[10221] = 8'h28;
mem[10222] = 8'h0e;
mem[10223] = 8'h03;
mem[10224] = 8'h02;
mem[10225] = 8'h08;
mem[10226] = 8'had;
mem[10227] = 8'h03;
mem[10228] = 8'h02;
mem[10229] = 8'hdd;
mem[10230] = 8'h20;
mem[10231] = 8'h02;
mem[10232] = 8'hd0;
mem[10233] = 8'hfe;
mem[10234] = 8'h68;
mem[10235] = 8'h09;
mem[10236] = 8'h08;
mem[10237] = 8'h49;
mem[10238] = 8'h38;
mem[10239] = 8'hdd;
mem[10240] = 8'h30;
mem[10241] = 8'h02;
mem[10242] = 8'hd0;
mem[10243] = 8'hfe;
mem[10244] = 8'hca;
mem[10245] = 8'h10;
mem[10246] = 8'hde;
mem[10247] = 8'ha2;
mem[10248] = 8'h03;
mem[10249] = 8'ha9;
mem[10250] = 8'hff;
mem[10251] = 8'h48;
mem[10252] = 8'hb5;
mem[10253] = 8'h13;
mem[10254] = 8'h8d;
mem[10255] = 8'h03;
mem[10256] = 8'h02;
mem[10257] = 8'h28;
mem[10258] = 8'h0e;
mem[10259] = 8'h03;
mem[10260] = 8'h02;
mem[10261] = 8'h08;
mem[10262] = 8'had;
mem[10263] = 8'h03;
mem[10264] = 8'h02;
mem[10265] = 8'hdd;
mem[10266] = 8'h20;
mem[10267] = 8'h02;
mem[10268] = 8'hd0;
mem[10269] = 8'hfe;
mem[10270] = 8'h68;
mem[10271] = 8'h09;
mem[10272] = 8'h08;
mem[10273] = 8'h49;
mem[10274] = 8'h7c;
mem[10275] = 8'hdd;
mem[10276] = 8'h30;
mem[10277] = 8'h02;
mem[10278] = 8'hd0;
mem[10279] = 8'hfe;
mem[10280] = 8'hca;
mem[10281] = 8'h10;
mem[10282] = 8'hde;
mem[10283] = 8'ha2;
mem[10284] = 8'h03;
mem[10285] = 8'ha9;
mem[10286] = 8'h00;
mem[10287] = 8'h48;
mem[10288] = 8'hb5;
mem[10289] = 8'h13;
mem[10290] = 8'h8d;
mem[10291] = 8'h03;
mem[10292] = 8'h02;
mem[10293] = 8'h28;
mem[10294] = 8'h4e;
mem[10295] = 8'h03;
mem[10296] = 8'h02;
mem[10297] = 8'h08;
mem[10298] = 8'had;
mem[10299] = 8'h03;
mem[10300] = 8'h02;
mem[10301] = 8'hdd;
mem[10302] = 8'h28;
mem[10303] = 8'h02;
mem[10304] = 8'hd0;
mem[10305] = 8'hfe;
mem[10306] = 8'h68;
mem[10307] = 8'h09;
mem[10308] = 8'h08;
mem[10309] = 8'h49;
mem[10310] = 8'h38;
mem[10311] = 8'hdd;
mem[10312] = 8'h38;
mem[10313] = 8'h02;
mem[10314] = 8'hd0;
mem[10315] = 8'hfe;
mem[10316] = 8'hca;
mem[10317] = 8'h10;
mem[10318] = 8'hde;
mem[10319] = 8'ha2;
mem[10320] = 8'h03;
mem[10321] = 8'ha9;
mem[10322] = 8'hff;
mem[10323] = 8'h48;
mem[10324] = 8'hb5;
mem[10325] = 8'h13;
mem[10326] = 8'h8d;
mem[10327] = 8'h03;
mem[10328] = 8'h02;
mem[10329] = 8'h28;
mem[10330] = 8'h4e;
mem[10331] = 8'h03;
mem[10332] = 8'h02;
mem[10333] = 8'h08;
mem[10334] = 8'had;
mem[10335] = 8'h03;
mem[10336] = 8'h02;
mem[10337] = 8'hdd;
mem[10338] = 8'h28;
mem[10339] = 8'h02;
mem[10340] = 8'hd0;
mem[10341] = 8'hfe;
mem[10342] = 8'h68;
mem[10343] = 8'h09;
mem[10344] = 8'h08;
mem[10345] = 8'h49;
mem[10346] = 8'h7c;
mem[10347] = 8'hdd;
mem[10348] = 8'h38;
mem[10349] = 8'h02;
mem[10350] = 8'hd0;
mem[10351] = 8'hfe;
mem[10352] = 8'hca;
mem[10353] = 8'h10;
mem[10354] = 8'hde;
mem[10355] = 8'ha2;
mem[10356] = 8'h03;
mem[10357] = 8'ha9;
mem[10358] = 8'h00;
mem[10359] = 8'h48;
mem[10360] = 8'hb5;
mem[10361] = 8'h13;
mem[10362] = 8'h8d;
mem[10363] = 8'h03;
mem[10364] = 8'h02;
mem[10365] = 8'h28;
mem[10366] = 8'h2e;
mem[10367] = 8'h03;
mem[10368] = 8'h02;
mem[10369] = 8'h08;
mem[10370] = 8'had;
mem[10371] = 8'h03;
mem[10372] = 8'h02;
mem[10373] = 8'hdd;
mem[10374] = 8'h20;
mem[10375] = 8'h02;
mem[10376] = 8'hd0;
mem[10377] = 8'hfe;
mem[10378] = 8'h68;
mem[10379] = 8'h09;
mem[10380] = 8'h08;
mem[10381] = 8'h49;
mem[10382] = 8'h38;
mem[10383] = 8'hdd;
mem[10384] = 8'h30;
mem[10385] = 8'h02;
mem[10386] = 8'hd0;
mem[10387] = 8'hfe;
mem[10388] = 8'hca;
mem[10389] = 8'h10;
mem[10390] = 8'hde;
mem[10391] = 8'ha2;
mem[10392] = 8'h03;
mem[10393] = 8'ha9;
mem[10394] = 8'hfe;
mem[10395] = 8'h48;
mem[10396] = 8'hb5;
mem[10397] = 8'h13;
mem[10398] = 8'h8d;
mem[10399] = 8'h03;
mem[10400] = 8'h02;
mem[10401] = 8'h28;
mem[10402] = 8'h2e;
mem[10403] = 8'h03;
mem[10404] = 8'h02;
mem[10405] = 8'h08;
mem[10406] = 8'had;
mem[10407] = 8'h03;
mem[10408] = 8'h02;
mem[10409] = 8'hdd;
mem[10410] = 8'h20;
mem[10411] = 8'h02;
mem[10412] = 8'hd0;
mem[10413] = 8'hfe;
mem[10414] = 8'h68;
mem[10415] = 8'h09;
mem[10416] = 8'h08;
mem[10417] = 8'h49;
mem[10418] = 8'h7c;
mem[10419] = 8'hdd;
mem[10420] = 8'h30;
mem[10421] = 8'h02;
mem[10422] = 8'hd0;
mem[10423] = 8'hfe;
mem[10424] = 8'hca;
mem[10425] = 8'h10;
mem[10426] = 8'hde;
mem[10427] = 8'ha2;
mem[10428] = 8'h03;
mem[10429] = 8'ha9;
mem[10430] = 8'h01;
mem[10431] = 8'h48;
mem[10432] = 8'hb5;
mem[10433] = 8'h13;
mem[10434] = 8'h8d;
mem[10435] = 8'h03;
mem[10436] = 8'h02;
mem[10437] = 8'h28;
mem[10438] = 8'h2e;
mem[10439] = 8'h03;
mem[10440] = 8'h02;
mem[10441] = 8'h08;
mem[10442] = 8'had;
mem[10443] = 8'h03;
mem[10444] = 8'h02;
mem[10445] = 8'hdd;
mem[10446] = 8'h24;
mem[10447] = 8'h02;
mem[10448] = 8'hd0;
mem[10449] = 8'hfe;
mem[10450] = 8'h68;
mem[10451] = 8'h09;
mem[10452] = 8'h08;
mem[10453] = 8'h49;
mem[10454] = 8'h38;
mem[10455] = 8'hdd;
mem[10456] = 8'h34;
mem[10457] = 8'h02;
mem[10458] = 8'hd0;
mem[10459] = 8'hfe;
mem[10460] = 8'hca;
mem[10461] = 8'h10;
mem[10462] = 8'hde;
mem[10463] = 8'ha2;
mem[10464] = 8'h03;
mem[10465] = 8'ha9;
mem[10466] = 8'hff;
mem[10467] = 8'h48;
mem[10468] = 8'hb5;
mem[10469] = 8'h13;
mem[10470] = 8'h8d;
mem[10471] = 8'h03;
mem[10472] = 8'h02;
mem[10473] = 8'h28;
mem[10474] = 8'h2e;
mem[10475] = 8'h03;
mem[10476] = 8'h02;
mem[10477] = 8'h08;
mem[10478] = 8'had;
mem[10479] = 8'h03;
mem[10480] = 8'h02;
mem[10481] = 8'hdd;
mem[10482] = 8'h24;
mem[10483] = 8'h02;
mem[10484] = 8'hd0;
mem[10485] = 8'hfe;
mem[10486] = 8'h68;
mem[10487] = 8'h09;
mem[10488] = 8'h08;
mem[10489] = 8'h49;
mem[10490] = 8'h7c;
mem[10491] = 8'hdd;
mem[10492] = 8'h34;
mem[10493] = 8'h02;
mem[10494] = 8'hd0;
mem[10495] = 8'hfe;
mem[10496] = 8'hca;
mem[10497] = 8'h10;
mem[10498] = 8'hde;
mem[10499] = 8'ha2;
mem[10500] = 8'h03;
mem[10501] = 8'ha9;
mem[10502] = 8'h00;
mem[10503] = 8'h48;
mem[10504] = 8'hb5;
mem[10505] = 8'h13;
mem[10506] = 8'h8d;
mem[10507] = 8'h03;
mem[10508] = 8'h02;
mem[10509] = 8'h28;
mem[10510] = 8'h6e;
mem[10511] = 8'h03;
mem[10512] = 8'h02;
mem[10513] = 8'h08;
mem[10514] = 8'had;
mem[10515] = 8'h03;
mem[10516] = 8'h02;
mem[10517] = 8'hdd;
mem[10518] = 8'h28;
mem[10519] = 8'h02;
mem[10520] = 8'hd0;
mem[10521] = 8'hfe;
mem[10522] = 8'h68;
mem[10523] = 8'h09;
mem[10524] = 8'h08;
mem[10525] = 8'h49;
mem[10526] = 8'h38;
mem[10527] = 8'hdd;
mem[10528] = 8'h38;
mem[10529] = 8'h02;
mem[10530] = 8'hd0;
mem[10531] = 8'hfe;
mem[10532] = 8'hca;
mem[10533] = 8'h10;
mem[10534] = 8'hde;
mem[10535] = 8'ha2;
mem[10536] = 8'h03;
mem[10537] = 8'ha9;
mem[10538] = 8'hfe;
mem[10539] = 8'h48;
mem[10540] = 8'hb5;
mem[10541] = 8'h13;
mem[10542] = 8'h8d;
mem[10543] = 8'h03;
mem[10544] = 8'h02;
mem[10545] = 8'h28;
mem[10546] = 8'h6e;
mem[10547] = 8'h03;
mem[10548] = 8'h02;
mem[10549] = 8'h08;
mem[10550] = 8'had;
mem[10551] = 8'h03;
mem[10552] = 8'h02;
mem[10553] = 8'hdd;
mem[10554] = 8'h28;
mem[10555] = 8'h02;
mem[10556] = 8'hd0;
mem[10557] = 8'hfe;
mem[10558] = 8'h68;
mem[10559] = 8'h09;
mem[10560] = 8'h08;
mem[10561] = 8'h49;
mem[10562] = 8'h7c;
mem[10563] = 8'hdd;
mem[10564] = 8'h38;
mem[10565] = 8'h02;
mem[10566] = 8'hd0;
mem[10567] = 8'hfe;
mem[10568] = 8'hca;
mem[10569] = 8'h10;
mem[10570] = 8'hde;
mem[10571] = 8'ha2;
mem[10572] = 8'h03;
mem[10573] = 8'ha9;
mem[10574] = 8'h01;
mem[10575] = 8'h48;
mem[10576] = 8'hb5;
mem[10577] = 8'h13;
mem[10578] = 8'h8d;
mem[10579] = 8'h03;
mem[10580] = 8'h02;
mem[10581] = 8'h28;
mem[10582] = 8'h6e;
mem[10583] = 8'h03;
mem[10584] = 8'h02;
mem[10585] = 8'h08;
mem[10586] = 8'had;
mem[10587] = 8'h03;
mem[10588] = 8'h02;
mem[10589] = 8'hdd;
mem[10590] = 8'h2c;
mem[10591] = 8'h02;
mem[10592] = 8'hd0;
mem[10593] = 8'hfe;
mem[10594] = 8'h68;
mem[10595] = 8'h09;
mem[10596] = 8'h08;
mem[10597] = 8'h49;
mem[10598] = 8'h38;
mem[10599] = 8'hdd;
mem[10600] = 8'h3c;
mem[10601] = 8'h02;
mem[10602] = 8'hd0;
mem[10603] = 8'hfe;
mem[10604] = 8'hca;
mem[10605] = 8'h10;
mem[10606] = 8'hde;
mem[10607] = 8'ha2;
mem[10608] = 8'h03;
mem[10609] = 8'ha9;
mem[10610] = 8'hff;
mem[10611] = 8'h48;
mem[10612] = 8'hb5;
mem[10613] = 8'h13;
mem[10614] = 8'h8d;
mem[10615] = 8'h03;
mem[10616] = 8'h02;
mem[10617] = 8'h28;
mem[10618] = 8'h6e;
mem[10619] = 8'h03;
mem[10620] = 8'h02;
mem[10621] = 8'h08;
mem[10622] = 8'had;
mem[10623] = 8'h03;
mem[10624] = 8'h02;
mem[10625] = 8'hdd;
mem[10626] = 8'h2c;
mem[10627] = 8'h02;
mem[10628] = 8'hd0;
mem[10629] = 8'hfe;
mem[10630] = 8'h68;
mem[10631] = 8'h09;
mem[10632] = 8'h08;
mem[10633] = 8'h49;
mem[10634] = 8'h7c;
mem[10635] = 8'hdd;
mem[10636] = 8'h3c;
mem[10637] = 8'h02;
mem[10638] = 8'hd0;
mem[10639] = 8'hfe;
mem[10640] = 8'hca;
mem[10641] = 8'h10;
mem[10642] = 8'hde;
mem[10643] = 8'had;
mem[10644] = 8'h00;
mem[10645] = 8'h02;
mem[10646] = 8'hc9;
mem[10647] = 8'h1f;
mem[10648] = 8'hd0;
mem[10649] = 8'hfe;
mem[10650] = 8'ha9;
mem[10651] = 8'h20;
mem[10652] = 8'h8d;
mem[10653] = 8'h00;
mem[10654] = 8'h02;
mem[10655] = 8'ha2;
mem[10656] = 8'h03;
mem[10657] = 8'ha9;
mem[10658] = 8'h00;
mem[10659] = 8'h48;
mem[10660] = 8'hb5;
mem[10661] = 8'h13;
mem[10662] = 8'h95;
mem[10663] = 8'h0c;
mem[10664] = 8'h28;
mem[10665] = 8'h16;
mem[10666] = 8'h0c;
mem[10667] = 8'h08;
mem[10668] = 8'hb5;
mem[10669] = 8'h0c;
mem[10670] = 8'hdd;
mem[10671] = 8'h20;
mem[10672] = 8'h02;
mem[10673] = 8'hd0;
mem[10674] = 8'hfe;
mem[10675] = 8'h68;
mem[10676] = 8'h09;
mem[10677] = 8'h08;
mem[10678] = 8'h49;
mem[10679] = 8'h38;
mem[10680] = 8'hdd;
mem[10681] = 8'h30;
mem[10682] = 8'h02;
mem[10683] = 8'hd0;
mem[10684] = 8'hfe;
mem[10685] = 8'hca;
mem[10686] = 8'h10;
mem[10687] = 8'he1;
mem[10688] = 8'ha2;
mem[10689] = 8'h03;
mem[10690] = 8'ha9;
mem[10691] = 8'hff;
mem[10692] = 8'h48;
mem[10693] = 8'hb5;
mem[10694] = 8'h13;
mem[10695] = 8'h95;
mem[10696] = 8'h0c;
mem[10697] = 8'h28;
mem[10698] = 8'h16;
mem[10699] = 8'h0c;
mem[10700] = 8'h08;
mem[10701] = 8'hb5;
mem[10702] = 8'h0c;
mem[10703] = 8'hdd;
mem[10704] = 8'h20;
mem[10705] = 8'h02;
mem[10706] = 8'hd0;
mem[10707] = 8'hfe;
mem[10708] = 8'h68;
mem[10709] = 8'h09;
mem[10710] = 8'h08;
mem[10711] = 8'h49;
mem[10712] = 8'h7c;
mem[10713] = 8'hdd;
mem[10714] = 8'h30;
mem[10715] = 8'h02;
mem[10716] = 8'hd0;
mem[10717] = 8'hfe;
mem[10718] = 8'hca;
mem[10719] = 8'h10;
mem[10720] = 8'he1;
mem[10721] = 8'ha2;
mem[10722] = 8'h03;
mem[10723] = 8'ha9;
mem[10724] = 8'h00;
mem[10725] = 8'h48;
mem[10726] = 8'hb5;
mem[10727] = 8'h13;
mem[10728] = 8'h95;
mem[10729] = 8'h0c;
mem[10730] = 8'h28;
mem[10731] = 8'h56;
mem[10732] = 8'h0c;
mem[10733] = 8'h08;
mem[10734] = 8'hb5;
mem[10735] = 8'h0c;
mem[10736] = 8'hdd;
mem[10737] = 8'h28;
mem[10738] = 8'h02;
mem[10739] = 8'hd0;
mem[10740] = 8'hfe;
mem[10741] = 8'h68;
mem[10742] = 8'h09;
mem[10743] = 8'h08;
mem[10744] = 8'h49;
mem[10745] = 8'h38;
mem[10746] = 8'hdd;
mem[10747] = 8'h38;
mem[10748] = 8'h02;
mem[10749] = 8'hd0;
mem[10750] = 8'hfe;
mem[10751] = 8'hca;
mem[10752] = 8'h10;
mem[10753] = 8'he1;
mem[10754] = 8'ha2;
mem[10755] = 8'h03;
mem[10756] = 8'ha9;
mem[10757] = 8'hff;
mem[10758] = 8'h48;
mem[10759] = 8'hb5;
mem[10760] = 8'h13;
mem[10761] = 8'h95;
mem[10762] = 8'h0c;
mem[10763] = 8'h28;
mem[10764] = 8'h56;
mem[10765] = 8'h0c;
mem[10766] = 8'h08;
mem[10767] = 8'hb5;
mem[10768] = 8'h0c;
mem[10769] = 8'hdd;
mem[10770] = 8'h28;
mem[10771] = 8'h02;
mem[10772] = 8'hd0;
mem[10773] = 8'hfe;
mem[10774] = 8'h68;
mem[10775] = 8'h09;
mem[10776] = 8'h08;
mem[10777] = 8'h49;
mem[10778] = 8'h7c;
mem[10779] = 8'hdd;
mem[10780] = 8'h38;
mem[10781] = 8'h02;
mem[10782] = 8'hd0;
mem[10783] = 8'hfe;
mem[10784] = 8'hca;
mem[10785] = 8'h10;
mem[10786] = 8'he1;
mem[10787] = 8'ha2;
mem[10788] = 8'h03;
mem[10789] = 8'ha9;
mem[10790] = 8'h00;
mem[10791] = 8'h48;
mem[10792] = 8'hb5;
mem[10793] = 8'h13;
mem[10794] = 8'h95;
mem[10795] = 8'h0c;
mem[10796] = 8'h28;
mem[10797] = 8'h36;
mem[10798] = 8'h0c;
mem[10799] = 8'h08;
mem[10800] = 8'hb5;
mem[10801] = 8'h0c;
mem[10802] = 8'hdd;
mem[10803] = 8'h20;
mem[10804] = 8'h02;
mem[10805] = 8'hd0;
mem[10806] = 8'hfe;
mem[10807] = 8'h68;
mem[10808] = 8'h09;
mem[10809] = 8'h08;
mem[10810] = 8'h49;
mem[10811] = 8'h38;
mem[10812] = 8'hdd;
mem[10813] = 8'h30;
mem[10814] = 8'h02;
mem[10815] = 8'hd0;
mem[10816] = 8'hfe;
mem[10817] = 8'hca;
mem[10818] = 8'h10;
mem[10819] = 8'he1;
mem[10820] = 8'ha2;
mem[10821] = 8'h03;
mem[10822] = 8'ha9;
mem[10823] = 8'hfe;
mem[10824] = 8'h48;
mem[10825] = 8'hb5;
mem[10826] = 8'h13;
mem[10827] = 8'h95;
mem[10828] = 8'h0c;
mem[10829] = 8'h28;
mem[10830] = 8'h36;
mem[10831] = 8'h0c;
mem[10832] = 8'h08;
mem[10833] = 8'hb5;
mem[10834] = 8'h0c;
mem[10835] = 8'hdd;
mem[10836] = 8'h20;
mem[10837] = 8'h02;
mem[10838] = 8'hd0;
mem[10839] = 8'hfe;
mem[10840] = 8'h68;
mem[10841] = 8'h09;
mem[10842] = 8'h08;
mem[10843] = 8'h49;
mem[10844] = 8'h7c;
mem[10845] = 8'hdd;
mem[10846] = 8'h30;
mem[10847] = 8'h02;
mem[10848] = 8'hd0;
mem[10849] = 8'hfe;
mem[10850] = 8'hca;
mem[10851] = 8'h10;
mem[10852] = 8'he1;
mem[10853] = 8'ha2;
mem[10854] = 8'h03;
mem[10855] = 8'ha9;
mem[10856] = 8'h01;
mem[10857] = 8'h48;
mem[10858] = 8'hb5;
mem[10859] = 8'h13;
mem[10860] = 8'h95;
mem[10861] = 8'h0c;
mem[10862] = 8'h28;
mem[10863] = 8'h36;
mem[10864] = 8'h0c;
mem[10865] = 8'h08;
mem[10866] = 8'hb5;
mem[10867] = 8'h0c;
mem[10868] = 8'hdd;
mem[10869] = 8'h24;
mem[10870] = 8'h02;
mem[10871] = 8'hd0;
mem[10872] = 8'hfe;
mem[10873] = 8'h68;
mem[10874] = 8'h09;
mem[10875] = 8'h08;
mem[10876] = 8'h49;
mem[10877] = 8'h38;
mem[10878] = 8'hdd;
mem[10879] = 8'h34;
mem[10880] = 8'h02;
mem[10881] = 8'hd0;
mem[10882] = 8'hfe;
mem[10883] = 8'hca;
mem[10884] = 8'h10;
mem[10885] = 8'he1;
mem[10886] = 8'ha2;
mem[10887] = 8'h03;
mem[10888] = 8'ha9;
mem[10889] = 8'hff;
mem[10890] = 8'h48;
mem[10891] = 8'hb5;
mem[10892] = 8'h13;
mem[10893] = 8'h95;
mem[10894] = 8'h0c;
mem[10895] = 8'h28;
mem[10896] = 8'h36;
mem[10897] = 8'h0c;
mem[10898] = 8'h08;
mem[10899] = 8'hb5;
mem[10900] = 8'h0c;
mem[10901] = 8'hdd;
mem[10902] = 8'h24;
mem[10903] = 8'h02;
mem[10904] = 8'hd0;
mem[10905] = 8'hfe;
mem[10906] = 8'h68;
mem[10907] = 8'h09;
mem[10908] = 8'h08;
mem[10909] = 8'h49;
mem[10910] = 8'h7c;
mem[10911] = 8'hdd;
mem[10912] = 8'h34;
mem[10913] = 8'h02;
mem[10914] = 8'hd0;
mem[10915] = 8'hfe;
mem[10916] = 8'hca;
mem[10917] = 8'h10;
mem[10918] = 8'he1;
mem[10919] = 8'ha2;
mem[10920] = 8'h03;
mem[10921] = 8'ha9;
mem[10922] = 8'h00;
mem[10923] = 8'h48;
mem[10924] = 8'hb5;
mem[10925] = 8'h13;
mem[10926] = 8'h95;
mem[10927] = 8'h0c;
mem[10928] = 8'h28;
mem[10929] = 8'h76;
mem[10930] = 8'h0c;
mem[10931] = 8'h08;
mem[10932] = 8'hb5;
mem[10933] = 8'h0c;
mem[10934] = 8'hdd;
mem[10935] = 8'h28;
mem[10936] = 8'h02;
mem[10937] = 8'hd0;
mem[10938] = 8'hfe;
mem[10939] = 8'h68;
mem[10940] = 8'h09;
mem[10941] = 8'h08;
mem[10942] = 8'h49;
mem[10943] = 8'h38;
mem[10944] = 8'hdd;
mem[10945] = 8'h38;
mem[10946] = 8'h02;
mem[10947] = 8'hd0;
mem[10948] = 8'hfe;
mem[10949] = 8'hca;
mem[10950] = 8'h10;
mem[10951] = 8'he1;
mem[10952] = 8'ha2;
mem[10953] = 8'h03;
mem[10954] = 8'ha9;
mem[10955] = 8'hfe;
mem[10956] = 8'h48;
mem[10957] = 8'hb5;
mem[10958] = 8'h13;
mem[10959] = 8'h95;
mem[10960] = 8'h0c;
mem[10961] = 8'h28;
mem[10962] = 8'h76;
mem[10963] = 8'h0c;
mem[10964] = 8'h08;
mem[10965] = 8'hb5;
mem[10966] = 8'h0c;
mem[10967] = 8'hdd;
mem[10968] = 8'h28;
mem[10969] = 8'h02;
mem[10970] = 8'hd0;
mem[10971] = 8'hfe;
mem[10972] = 8'h68;
mem[10973] = 8'h09;
mem[10974] = 8'h08;
mem[10975] = 8'h49;
mem[10976] = 8'h7c;
mem[10977] = 8'hdd;
mem[10978] = 8'h38;
mem[10979] = 8'h02;
mem[10980] = 8'hd0;
mem[10981] = 8'hfe;
mem[10982] = 8'hca;
mem[10983] = 8'h10;
mem[10984] = 8'he1;
mem[10985] = 8'ha2;
mem[10986] = 8'h03;
mem[10987] = 8'ha9;
mem[10988] = 8'h01;
mem[10989] = 8'h48;
mem[10990] = 8'hb5;
mem[10991] = 8'h13;
mem[10992] = 8'h95;
mem[10993] = 8'h0c;
mem[10994] = 8'h28;
mem[10995] = 8'h76;
mem[10996] = 8'h0c;
mem[10997] = 8'h08;
mem[10998] = 8'hb5;
mem[10999] = 8'h0c;
mem[11000] = 8'hdd;
mem[11001] = 8'h2c;
mem[11002] = 8'h02;
mem[11003] = 8'hd0;
mem[11004] = 8'hfe;
mem[11005] = 8'h68;
mem[11006] = 8'h09;
mem[11007] = 8'h08;
mem[11008] = 8'h49;
mem[11009] = 8'h38;
mem[11010] = 8'hdd;
mem[11011] = 8'h3c;
mem[11012] = 8'h02;
mem[11013] = 8'hd0;
mem[11014] = 8'hfe;
mem[11015] = 8'hca;
mem[11016] = 8'h10;
mem[11017] = 8'he1;
mem[11018] = 8'ha2;
mem[11019] = 8'h03;
mem[11020] = 8'ha9;
mem[11021] = 8'hff;
mem[11022] = 8'h48;
mem[11023] = 8'hb5;
mem[11024] = 8'h13;
mem[11025] = 8'h95;
mem[11026] = 8'h0c;
mem[11027] = 8'h28;
mem[11028] = 8'h76;
mem[11029] = 8'h0c;
mem[11030] = 8'h08;
mem[11031] = 8'hb5;
mem[11032] = 8'h0c;
mem[11033] = 8'hdd;
mem[11034] = 8'h2c;
mem[11035] = 8'h02;
mem[11036] = 8'hd0;
mem[11037] = 8'hfe;
mem[11038] = 8'h68;
mem[11039] = 8'h09;
mem[11040] = 8'h08;
mem[11041] = 8'h49;
mem[11042] = 8'h7c;
mem[11043] = 8'hdd;
mem[11044] = 8'h3c;
mem[11045] = 8'h02;
mem[11046] = 8'hd0;
mem[11047] = 8'hfe;
mem[11048] = 8'hca;
mem[11049] = 8'h10;
mem[11050] = 8'he1;
mem[11051] = 8'had;
mem[11052] = 8'h00;
mem[11053] = 8'h02;
mem[11054] = 8'hc9;
mem[11055] = 8'h20;
mem[11056] = 8'hd0;
mem[11057] = 8'hfe;
mem[11058] = 8'ha9;
mem[11059] = 8'h21;
mem[11060] = 8'h8d;
mem[11061] = 8'h00;
mem[11062] = 8'h02;
mem[11063] = 8'ha2;
mem[11064] = 8'h03;
mem[11065] = 8'ha9;
mem[11066] = 8'h00;
mem[11067] = 8'h48;
mem[11068] = 8'hb5;
mem[11069] = 8'h13;
mem[11070] = 8'h9d;
mem[11071] = 8'h03;
mem[11072] = 8'h02;
mem[11073] = 8'h28;
mem[11074] = 8'h1e;
mem[11075] = 8'h03;
mem[11076] = 8'h02;
mem[11077] = 8'h08;
mem[11078] = 8'hbd;
mem[11079] = 8'h03;
mem[11080] = 8'h02;
mem[11081] = 8'hdd;
mem[11082] = 8'h20;
mem[11083] = 8'h02;
mem[11084] = 8'hd0;
mem[11085] = 8'hfe;
mem[11086] = 8'h68;
mem[11087] = 8'h09;
mem[11088] = 8'h08;
mem[11089] = 8'h49;
mem[11090] = 8'h38;
mem[11091] = 8'hdd;
mem[11092] = 8'h30;
mem[11093] = 8'h02;
mem[11094] = 8'hd0;
mem[11095] = 8'hfe;
mem[11096] = 8'hca;
mem[11097] = 8'h10;
mem[11098] = 8'hde;
mem[11099] = 8'ha2;
mem[11100] = 8'h03;
mem[11101] = 8'ha9;
mem[11102] = 8'hff;
mem[11103] = 8'h48;
mem[11104] = 8'hb5;
mem[11105] = 8'h13;
mem[11106] = 8'h9d;
mem[11107] = 8'h03;
mem[11108] = 8'h02;
mem[11109] = 8'h28;
mem[11110] = 8'h1e;
mem[11111] = 8'h03;
mem[11112] = 8'h02;
mem[11113] = 8'h08;
mem[11114] = 8'hbd;
mem[11115] = 8'h03;
mem[11116] = 8'h02;
mem[11117] = 8'hdd;
mem[11118] = 8'h20;
mem[11119] = 8'h02;
mem[11120] = 8'hd0;
mem[11121] = 8'hfe;
mem[11122] = 8'h68;
mem[11123] = 8'h09;
mem[11124] = 8'h08;
mem[11125] = 8'h49;
mem[11126] = 8'h7c;
mem[11127] = 8'hdd;
mem[11128] = 8'h30;
mem[11129] = 8'h02;
mem[11130] = 8'hd0;
mem[11131] = 8'hfe;
mem[11132] = 8'hca;
mem[11133] = 8'h10;
mem[11134] = 8'hde;
mem[11135] = 8'ha2;
mem[11136] = 8'h03;
mem[11137] = 8'ha9;
mem[11138] = 8'h00;
mem[11139] = 8'h48;
mem[11140] = 8'hb5;
mem[11141] = 8'h13;
mem[11142] = 8'h9d;
mem[11143] = 8'h03;
mem[11144] = 8'h02;
mem[11145] = 8'h28;
mem[11146] = 8'h5e;
mem[11147] = 8'h03;
mem[11148] = 8'h02;
mem[11149] = 8'h08;
mem[11150] = 8'hbd;
mem[11151] = 8'h03;
mem[11152] = 8'h02;
mem[11153] = 8'hdd;
mem[11154] = 8'h28;
mem[11155] = 8'h02;
mem[11156] = 8'hd0;
mem[11157] = 8'hfe;
mem[11158] = 8'h68;
mem[11159] = 8'h09;
mem[11160] = 8'h08;
mem[11161] = 8'h49;
mem[11162] = 8'h38;
mem[11163] = 8'hdd;
mem[11164] = 8'h38;
mem[11165] = 8'h02;
mem[11166] = 8'hd0;
mem[11167] = 8'hfe;
mem[11168] = 8'hca;
mem[11169] = 8'h10;
mem[11170] = 8'hde;
mem[11171] = 8'ha2;
mem[11172] = 8'h03;
mem[11173] = 8'ha9;
mem[11174] = 8'hff;
mem[11175] = 8'h48;
mem[11176] = 8'hb5;
mem[11177] = 8'h13;
mem[11178] = 8'h9d;
mem[11179] = 8'h03;
mem[11180] = 8'h02;
mem[11181] = 8'h28;
mem[11182] = 8'h5e;
mem[11183] = 8'h03;
mem[11184] = 8'h02;
mem[11185] = 8'h08;
mem[11186] = 8'hbd;
mem[11187] = 8'h03;
mem[11188] = 8'h02;
mem[11189] = 8'hdd;
mem[11190] = 8'h28;
mem[11191] = 8'h02;
mem[11192] = 8'hd0;
mem[11193] = 8'hfe;
mem[11194] = 8'h68;
mem[11195] = 8'h09;
mem[11196] = 8'h08;
mem[11197] = 8'h49;
mem[11198] = 8'h7c;
mem[11199] = 8'hdd;
mem[11200] = 8'h38;
mem[11201] = 8'h02;
mem[11202] = 8'hd0;
mem[11203] = 8'hfe;
mem[11204] = 8'hca;
mem[11205] = 8'h10;
mem[11206] = 8'hde;
mem[11207] = 8'ha2;
mem[11208] = 8'h03;
mem[11209] = 8'ha9;
mem[11210] = 8'h00;
mem[11211] = 8'h48;
mem[11212] = 8'hb5;
mem[11213] = 8'h13;
mem[11214] = 8'h9d;
mem[11215] = 8'h03;
mem[11216] = 8'h02;
mem[11217] = 8'h28;
mem[11218] = 8'h3e;
mem[11219] = 8'h03;
mem[11220] = 8'h02;
mem[11221] = 8'h08;
mem[11222] = 8'hbd;
mem[11223] = 8'h03;
mem[11224] = 8'h02;
mem[11225] = 8'hdd;
mem[11226] = 8'h20;
mem[11227] = 8'h02;
mem[11228] = 8'hd0;
mem[11229] = 8'hfe;
mem[11230] = 8'h68;
mem[11231] = 8'h09;
mem[11232] = 8'h08;
mem[11233] = 8'h49;
mem[11234] = 8'h38;
mem[11235] = 8'hdd;
mem[11236] = 8'h30;
mem[11237] = 8'h02;
mem[11238] = 8'hd0;
mem[11239] = 8'hfe;
mem[11240] = 8'hca;
mem[11241] = 8'h10;
mem[11242] = 8'hde;
mem[11243] = 8'ha2;
mem[11244] = 8'h03;
mem[11245] = 8'ha9;
mem[11246] = 8'hfe;
mem[11247] = 8'h48;
mem[11248] = 8'hb5;
mem[11249] = 8'h13;
mem[11250] = 8'h9d;
mem[11251] = 8'h03;
mem[11252] = 8'h02;
mem[11253] = 8'h28;
mem[11254] = 8'h3e;
mem[11255] = 8'h03;
mem[11256] = 8'h02;
mem[11257] = 8'h08;
mem[11258] = 8'hbd;
mem[11259] = 8'h03;
mem[11260] = 8'h02;
mem[11261] = 8'hdd;
mem[11262] = 8'h20;
mem[11263] = 8'h02;
mem[11264] = 8'hd0;
mem[11265] = 8'hfe;
mem[11266] = 8'h68;
mem[11267] = 8'h09;
mem[11268] = 8'h08;
mem[11269] = 8'h49;
mem[11270] = 8'h7c;
mem[11271] = 8'hdd;
mem[11272] = 8'h30;
mem[11273] = 8'h02;
mem[11274] = 8'hd0;
mem[11275] = 8'hfe;
mem[11276] = 8'hca;
mem[11277] = 8'h10;
mem[11278] = 8'hde;
mem[11279] = 8'ha2;
mem[11280] = 8'h03;
mem[11281] = 8'ha9;
mem[11282] = 8'h01;
mem[11283] = 8'h48;
mem[11284] = 8'hb5;
mem[11285] = 8'h13;
mem[11286] = 8'h9d;
mem[11287] = 8'h03;
mem[11288] = 8'h02;
mem[11289] = 8'h28;
mem[11290] = 8'h3e;
mem[11291] = 8'h03;
mem[11292] = 8'h02;
mem[11293] = 8'h08;
mem[11294] = 8'hbd;
mem[11295] = 8'h03;
mem[11296] = 8'h02;
mem[11297] = 8'hdd;
mem[11298] = 8'h24;
mem[11299] = 8'h02;
mem[11300] = 8'hd0;
mem[11301] = 8'hfe;
mem[11302] = 8'h68;
mem[11303] = 8'h09;
mem[11304] = 8'h08;
mem[11305] = 8'h49;
mem[11306] = 8'h38;
mem[11307] = 8'hdd;
mem[11308] = 8'h34;
mem[11309] = 8'h02;
mem[11310] = 8'hd0;
mem[11311] = 8'hfe;
mem[11312] = 8'hca;
mem[11313] = 8'h10;
mem[11314] = 8'hde;
mem[11315] = 8'ha2;
mem[11316] = 8'h03;
mem[11317] = 8'ha9;
mem[11318] = 8'hff;
mem[11319] = 8'h48;
mem[11320] = 8'hb5;
mem[11321] = 8'h13;
mem[11322] = 8'h9d;
mem[11323] = 8'h03;
mem[11324] = 8'h02;
mem[11325] = 8'h28;
mem[11326] = 8'h3e;
mem[11327] = 8'h03;
mem[11328] = 8'h02;
mem[11329] = 8'h08;
mem[11330] = 8'hbd;
mem[11331] = 8'h03;
mem[11332] = 8'h02;
mem[11333] = 8'hdd;
mem[11334] = 8'h24;
mem[11335] = 8'h02;
mem[11336] = 8'hd0;
mem[11337] = 8'hfe;
mem[11338] = 8'h68;
mem[11339] = 8'h09;
mem[11340] = 8'h08;
mem[11341] = 8'h49;
mem[11342] = 8'h7c;
mem[11343] = 8'hdd;
mem[11344] = 8'h34;
mem[11345] = 8'h02;
mem[11346] = 8'hd0;
mem[11347] = 8'hfe;
mem[11348] = 8'hca;
mem[11349] = 8'h10;
mem[11350] = 8'hde;
mem[11351] = 8'ha2;
mem[11352] = 8'h03;
mem[11353] = 8'ha9;
mem[11354] = 8'h00;
mem[11355] = 8'h48;
mem[11356] = 8'hb5;
mem[11357] = 8'h13;
mem[11358] = 8'h9d;
mem[11359] = 8'h03;
mem[11360] = 8'h02;
mem[11361] = 8'h28;
mem[11362] = 8'h7e;
mem[11363] = 8'h03;
mem[11364] = 8'h02;
mem[11365] = 8'h08;
mem[11366] = 8'hbd;
mem[11367] = 8'h03;
mem[11368] = 8'h02;
mem[11369] = 8'hdd;
mem[11370] = 8'h28;
mem[11371] = 8'h02;
mem[11372] = 8'hd0;
mem[11373] = 8'hfe;
mem[11374] = 8'h68;
mem[11375] = 8'h09;
mem[11376] = 8'h08;
mem[11377] = 8'h49;
mem[11378] = 8'h38;
mem[11379] = 8'hdd;
mem[11380] = 8'h38;
mem[11381] = 8'h02;
mem[11382] = 8'hd0;
mem[11383] = 8'hfe;
mem[11384] = 8'hca;
mem[11385] = 8'h10;
mem[11386] = 8'hde;
mem[11387] = 8'ha2;
mem[11388] = 8'h03;
mem[11389] = 8'ha9;
mem[11390] = 8'hfe;
mem[11391] = 8'h48;
mem[11392] = 8'hb5;
mem[11393] = 8'h13;
mem[11394] = 8'h9d;
mem[11395] = 8'h03;
mem[11396] = 8'h02;
mem[11397] = 8'h28;
mem[11398] = 8'h7e;
mem[11399] = 8'h03;
mem[11400] = 8'h02;
mem[11401] = 8'h08;
mem[11402] = 8'hbd;
mem[11403] = 8'h03;
mem[11404] = 8'h02;
mem[11405] = 8'hdd;
mem[11406] = 8'h28;
mem[11407] = 8'h02;
mem[11408] = 8'hd0;
mem[11409] = 8'hfe;
mem[11410] = 8'h68;
mem[11411] = 8'h09;
mem[11412] = 8'h08;
mem[11413] = 8'h49;
mem[11414] = 8'h7c;
mem[11415] = 8'hdd;
mem[11416] = 8'h38;
mem[11417] = 8'h02;
mem[11418] = 8'hd0;
mem[11419] = 8'hfe;
mem[11420] = 8'hca;
mem[11421] = 8'h10;
mem[11422] = 8'hde;
mem[11423] = 8'ha2;
mem[11424] = 8'h03;
mem[11425] = 8'ha9;
mem[11426] = 8'h01;
mem[11427] = 8'h48;
mem[11428] = 8'hb5;
mem[11429] = 8'h13;
mem[11430] = 8'h9d;
mem[11431] = 8'h03;
mem[11432] = 8'h02;
mem[11433] = 8'h28;
mem[11434] = 8'h7e;
mem[11435] = 8'h03;
mem[11436] = 8'h02;
mem[11437] = 8'h08;
mem[11438] = 8'hbd;
mem[11439] = 8'h03;
mem[11440] = 8'h02;
mem[11441] = 8'hdd;
mem[11442] = 8'h2c;
mem[11443] = 8'h02;
mem[11444] = 8'hd0;
mem[11445] = 8'hfe;
mem[11446] = 8'h68;
mem[11447] = 8'h09;
mem[11448] = 8'h08;
mem[11449] = 8'h49;
mem[11450] = 8'h38;
mem[11451] = 8'hdd;
mem[11452] = 8'h3c;
mem[11453] = 8'h02;
mem[11454] = 8'hd0;
mem[11455] = 8'hfe;
mem[11456] = 8'hca;
mem[11457] = 8'h10;
mem[11458] = 8'hde;
mem[11459] = 8'ha2;
mem[11460] = 8'h03;
mem[11461] = 8'ha9;
mem[11462] = 8'hff;
mem[11463] = 8'h48;
mem[11464] = 8'hb5;
mem[11465] = 8'h13;
mem[11466] = 8'h9d;
mem[11467] = 8'h03;
mem[11468] = 8'h02;
mem[11469] = 8'h28;
mem[11470] = 8'h7e;
mem[11471] = 8'h03;
mem[11472] = 8'h02;
mem[11473] = 8'h08;
mem[11474] = 8'hbd;
mem[11475] = 8'h03;
mem[11476] = 8'h02;
mem[11477] = 8'hdd;
mem[11478] = 8'h2c;
mem[11479] = 8'h02;
mem[11480] = 8'hd0;
mem[11481] = 8'hfe;
mem[11482] = 8'h68;
mem[11483] = 8'h09;
mem[11484] = 8'h08;
mem[11485] = 8'h49;
mem[11486] = 8'h7c;
mem[11487] = 8'hdd;
mem[11488] = 8'h3c;
mem[11489] = 8'h02;
mem[11490] = 8'hd0;
mem[11491] = 8'hfe;
mem[11492] = 8'hca;
mem[11493] = 8'h10;
mem[11494] = 8'hde;
mem[11495] = 8'had;
mem[11496] = 8'h00;
mem[11497] = 8'h02;
mem[11498] = 8'hc9;
mem[11499] = 8'h21;
mem[11500] = 8'hd0;
mem[11501] = 8'hfe;
mem[11502] = 8'ha9;
mem[11503] = 8'h22;
mem[11504] = 8'h8d;
mem[11505] = 8'h00;
mem[11506] = 8'h02;
mem[11507] = 8'ha2;
mem[11508] = 8'h00;
mem[11509] = 8'ha9;
mem[11510] = 8'h7e;
mem[11511] = 8'h85;
mem[11512] = 8'h0c;
mem[11513] = 8'ha9;
mem[11514] = 8'h00;
mem[11515] = 8'h48;
mem[11516] = 8'h28;
mem[11517] = 8'he6;
mem[11518] = 8'h0c;
mem[11519] = 8'h08;
mem[11520] = 8'ha5;
mem[11521] = 8'h0c;
mem[11522] = 8'hdd;
mem[11523] = 8'h40;
mem[11524] = 8'h02;
mem[11525] = 8'hd0;
mem[11526] = 8'hfe;
mem[11527] = 8'h68;
mem[11528] = 8'h09;
mem[11529] = 8'h08;
mem[11530] = 8'h49;
mem[11531] = 8'h38;
mem[11532] = 8'hdd;
mem[11533] = 8'h45;
mem[11534] = 8'h02;
mem[11535] = 8'hd0;
mem[11536] = 8'hfe;
mem[11537] = 8'he8;
mem[11538] = 8'he0;
mem[11539] = 8'h02;
mem[11540] = 8'hd0;
mem[11541] = 8'h04;
mem[11542] = 8'ha9;
mem[11543] = 8'hfe;
mem[11544] = 8'h85;
mem[11545] = 8'h0c;
mem[11546] = 8'he0;
mem[11547] = 8'h05;
mem[11548] = 8'hd0;
mem[11549] = 8'hdb;
mem[11550] = 8'hca;
mem[11551] = 8'he6;
mem[11552] = 8'h0c;
mem[11553] = 8'ha9;
mem[11554] = 8'h00;
mem[11555] = 8'h48;
mem[11556] = 8'h28;
mem[11557] = 8'hc6;
mem[11558] = 8'h0c;
mem[11559] = 8'h08;
mem[11560] = 8'ha5;
mem[11561] = 8'h0c;
mem[11562] = 8'hdd;
mem[11563] = 8'h40;
mem[11564] = 8'h02;
mem[11565] = 8'hd0;
mem[11566] = 8'hfe;
mem[11567] = 8'h68;
mem[11568] = 8'h09;
mem[11569] = 8'h08;
mem[11570] = 8'h49;
mem[11571] = 8'h38;
mem[11572] = 8'hdd;
mem[11573] = 8'h45;
mem[11574] = 8'h02;
mem[11575] = 8'hd0;
mem[11576] = 8'hfe;
mem[11577] = 8'hca;
mem[11578] = 8'h30;
mem[11579] = 8'h0a;
mem[11580] = 8'he0;
mem[11581] = 8'h01;
mem[11582] = 8'hd0;
mem[11583] = 8'he1;
mem[11584] = 8'ha9;
mem[11585] = 8'h81;
mem[11586] = 8'h85;
mem[11587] = 8'h0c;
mem[11588] = 8'hd0;
mem[11589] = 8'hdb;
mem[11590] = 8'ha2;
mem[11591] = 8'h00;
mem[11592] = 8'ha9;
mem[11593] = 8'h7e;
mem[11594] = 8'h85;
mem[11595] = 8'h0c;
mem[11596] = 8'ha9;
mem[11597] = 8'hff;
mem[11598] = 8'h48;
mem[11599] = 8'h28;
mem[11600] = 8'he6;
mem[11601] = 8'h0c;
mem[11602] = 8'h08;
mem[11603] = 8'ha5;
mem[11604] = 8'h0c;
mem[11605] = 8'hdd;
mem[11606] = 8'h40;
mem[11607] = 8'h02;
mem[11608] = 8'hd0;
mem[11609] = 8'hfe;
mem[11610] = 8'h68;
mem[11611] = 8'h09;
mem[11612] = 8'h08;
mem[11613] = 8'h49;
mem[11614] = 8'h7d;
mem[11615] = 8'hdd;
mem[11616] = 8'h45;
mem[11617] = 8'h02;
mem[11618] = 8'hd0;
mem[11619] = 8'hfe;
mem[11620] = 8'he8;
mem[11621] = 8'he0;
mem[11622] = 8'h02;
mem[11623] = 8'hd0;
mem[11624] = 8'h04;
mem[11625] = 8'ha9;
mem[11626] = 8'hfe;
mem[11627] = 8'h85;
mem[11628] = 8'h0c;
mem[11629] = 8'he0;
mem[11630] = 8'h05;
mem[11631] = 8'hd0;
mem[11632] = 8'hdb;
mem[11633] = 8'hca;
mem[11634] = 8'he6;
mem[11635] = 8'h0c;
mem[11636] = 8'ha9;
mem[11637] = 8'hff;
mem[11638] = 8'h48;
mem[11639] = 8'h28;
mem[11640] = 8'hc6;
mem[11641] = 8'h0c;
mem[11642] = 8'h08;
mem[11643] = 8'ha5;
mem[11644] = 8'h0c;
mem[11645] = 8'hdd;
mem[11646] = 8'h40;
mem[11647] = 8'h02;
mem[11648] = 8'hd0;
mem[11649] = 8'hfe;
mem[11650] = 8'h68;
mem[11651] = 8'h09;
mem[11652] = 8'h08;
mem[11653] = 8'h49;
mem[11654] = 8'h7d;
mem[11655] = 8'hdd;
mem[11656] = 8'h45;
mem[11657] = 8'h02;
mem[11658] = 8'hd0;
mem[11659] = 8'hfe;
mem[11660] = 8'hca;
mem[11661] = 8'h30;
mem[11662] = 8'h0a;
mem[11663] = 8'he0;
mem[11664] = 8'h01;
mem[11665] = 8'hd0;
mem[11666] = 8'he1;
mem[11667] = 8'ha9;
mem[11668] = 8'h81;
mem[11669] = 8'h85;
mem[11670] = 8'h0c;
mem[11671] = 8'hd0;
mem[11672] = 8'hdb;
mem[11673] = 8'had;
mem[11674] = 8'h00;
mem[11675] = 8'h02;
mem[11676] = 8'hc9;
mem[11677] = 8'h22;
mem[11678] = 8'hd0;
mem[11679] = 8'hfe;
mem[11680] = 8'ha9;
mem[11681] = 8'h23;
mem[11682] = 8'h8d;
mem[11683] = 8'h00;
mem[11684] = 8'h02;
mem[11685] = 8'ha2;
mem[11686] = 8'h00;
mem[11687] = 8'ha9;
mem[11688] = 8'h7e;
mem[11689] = 8'h8d;
mem[11690] = 8'h03;
mem[11691] = 8'h02;
mem[11692] = 8'ha9;
mem[11693] = 8'h00;
mem[11694] = 8'h48;
mem[11695] = 8'h28;
mem[11696] = 8'hee;
mem[11697] = 8'h03;
mem[11698] = 8'h02;
mem[11699] = 8'h08;
mem[11700] = 8'had;
mem[11701] = 8'h03;
mem[11702] = 8'h02;
mem[11703] = 8'hdd;
mem[11704] = 8'h40;
mem[11705] = 8'h02;
mem[11706] = 8'hd0;
mem[11707] = 8'hfe;
mem[11708] = 8'h68;
mem[11709] = 8'h09;
mem[11710] = 8'h08;
mem[11711] = 8'h49;
mem[11712] = 8'h38;
mem[11713] = 8'hdd;
mem[11714] = 8'h45;
mem[11715] = 8'h02;
mem[11716] = 8'hd0;
mem[11717] = 8'hfe;
mem[11718] = 8'he8;
mem[11719] = 8'he0;
mem[11720] = 8'h02;
mem[11721] = 8'hd0;
mem[11722] = 8'h05;
mem[11723] = 8'ha9;
mem[11724] = 8'hfe;
mem[11725] = 8'h8d;
mem[11726] = 8'h03;
mem[11727] = 8'h02;
mem[11728] = 8'he0;
mem[11729] = 8'h05;
mem[11730] = 8'hd0;
mem[11731] = 8'hd8;
mem[11732] = 8'hca;
mem[11733] = 8'hee;
mem[11734] = 8'h03;
mem[11735] = 8'h02;
mem[11736] = 8'ha9;
mem[11737] = 8'h00;
mem[11738] = 8'h48;
mem[11739] = 8'h28;
mem[11740] = 8'hce;
mem[11741] = 8'h03;
mem[11742] = 8'h02;
mem[11743] = 8'h08;
mem[11744] = 8'had;
mem[11745] = 8'h03;
mem[11746] = 8'h02;
mem[11747] = 8'hdd;
mem[11748] = 8'h40;
mem[11749] = 8'h02;
mem[11750] = 8'hd0;
mem[11751] = 8'hfe;
mem[11752] = 8'h68;
mem[11753] = 8'h09;
mem[11754] = 8'h08;
mem[11755] = 8'h49;
mem[11756] = 8'h38;
mem[11757] = 8'hdd;
mem[11758] = 8'h45;
mem[11759] = 8'h02;
mem[11760] = 8'hd0;
mem[11761] = 8'hfe;
mem[11762] = 8'hca;
mem[11763] = 8'h30;
mem[11764] = 8'h0b;
mem[11765] = 8'he0;
mem[11766] = 8'h01;
mem[11767] = 8'hd0;
mem[11768] = 8'hdf;
mem[11769] = 8'ha9;
mem[11770] = 8'h81;
mem[11771] = 8'h8d;
mem[11772] = 8'h03;
mem[11773] = 8'h02;
mem[11774] = 8'hd0;
mem[11775] = 8'hd8;
mem[11776] = 8'ha2;
mem[11777] = 8'h00;
mem[11778] = 8'ha9;
mem[11779] = 8'h7e;
mem[11780] = 8'h8d;
mem[11781] = 8'h03;
mem[11782] = 8'h02;
mem[11783] = 8'ha9;
mem[11784] = 8'hff;
mem[11785] = 8'h48;
mem[11786] = 8'h28;
mem[11787] = 8'hee;
mem[11788] = 8'h03;
mem[11789] = 8'h02;
mem[11790] = 8'h08;
mem[11791] = 8'had;
mem[11792] = 8'h03;
mem[11793] = 8'h02;
mem[11794] = 8'hdd;
mem[11795] = 8'h40;
mem[11796] = 8'h02;
mem[11797] = 8'hd0;
mem[11798] = 8'hfe;
mem[11799] = 8'h68;
mem[11800] = 8'h09;
mem[11801] = 8'h08;
mem[11802] = 8'h49;
mem[11803] = 8'h7d;
mem[11804] = 8'hdd;
mem[11805] = 8'h45;
mem[11806] = 8'h02;
mem[11807] = 8'hd0;
mem[11808] = 8'hfe;
mem[11809] = 8'he8;
mem[11810] = 8'he0;
mem[11811] = 8'h02;
mem[11812] = 8'hd0;
mem[11813] = 8'h05;
mem[11814] = 8'ha9;
mem[11815] = 8'hfe;
mem[11816] = 8'h8d;
mem[11817] = 8'h03;
mem[11818] = 8'h02;
mem[11819] = 8'he0;
mem[11820] = 8'h05;
mem[11821] = 8'hd0;
mem[11822] = 8'hd8;
mem[11823] = 8'hca;
mem[11824] = 8'hee;
mem[11825] = 8'h03;
mem[11826] = 8'h02;
mem[11827] = 8'ha9;
mem[11828] = 8'hff;
mem[11829] = 8'h48;
mem[11830] = 8'h28;
mem[11831] = 8'hce;
mem[11832] = 8'h03;
mem[11833] = 8'h02;
mem[11834] = 8'h08;
mem[11835] = 8'had;
mem[11836] = 8'h03;
mem[11837] = 8'h02;
mem[11838] = 8'hdd;
mem[11839] = 8'h40;
mem[11840] = 8'h02;
mem[11841] = 8'hd0;
mem[11842] = 8'hfe;
mem[11843] = 8'h68;
mem[11844] = 8'h09;
mem[11845] = 8'h08;
mem[11846] = 8'h49;
mem[11847] = 8'h7d;
mem[11848] = 8'hdd;
mem[11849] = 8'h45;
mem[11850] = 8'h02;
mem[11851] = 8'hd0;
mem[11852] = 8'hfe;
mem[11853] = 8'hca;
mem[11854] = 8'h30;
mem[11855] = 8'h0b;
mem[11856] = 8'he0;
mem[11857] = 8'h01;
mem[11858] = 8'hd0;
mem[11859] = 8'hdf;
mem[11860] = 8'ha9;
mem[11861] = 8'h81;
mem[11862] = 8'h8d;
mem[11863] = 8'h03;
mem[11864] = 8'h02;
mem[11865] = 8'hd0;
mem[11866] = 8'hd8;
mem[11867] = 8'had;
mem[11868] = 8'h00;
mem[11869] = 8'h02;
mem[11870] = 8'hc9;
mem[11871] = 8'h23;
mem[11872] = 8'hd0;
mem[11873] = 8'hfe;
mem[11874] = 8'ha9;
mem[11875] = 8'h24;
mem[11876] = 8'h8d;
mem[11877] = 8'h00;
mem[11878] = 8'h02;
mem[11879] = 8'ha2;
mem[11880] = 8'h00;
mem[11881] = 8'ha9;
mem[11882] = 8'h7e;
mem[11883] = 8'h95;
mem[11884] = 8'h0c;
mem[11885] = 8'ha9;
mem[11886] = 8'h00;
mem[11887] = 8'h48;
mem[11888] = 8'h28;
mem[11889] = 8'hf6;
mem[11890] = 8'h0c;
mem[11891] = 8'h08;
mem[11892] = 8'hb5;
mem[11893] = 8'h0c;
mem[11894] = 8'hdd;
mem[11895] = 8'h40;
mem[11896] = 8'h02;
mem[11897] = 8'hd0;
mem[11898] = 8'hfe;
mem[11899] = 8'h68;
mem[11900] = 8'h09;
mem[11901] = 8'h08;
mem[11902] = 8'h49;
mem[11903] = 8'h38;
mem[11904] = 8'hdd;
mem[11905] = 8'h45;
mem[11906] = 8'h02;
mem[11907] = 8'hd0;
mem[11908] = 8'hfe;
mem[11909] = 8'hb5;
mem[11910] = 8'h0c;
mem[11911] = 8'he8;
mem[11912] = 8'he0;
mem[11913] = 8'h02;
mem[11914] = 8'hd0;
mem[11915] = 8'h02;
mem[11916] = 8'ha9;
mem[11917] = 8'hfe;
mem[11918] = 8'he0;
mem[11919] = 8'h05;
mem[11920] = 8'hd0;
mem[11921] = 8'hd9;
mem[11922] = 8'hca;
mem[11923] = 8'ha9;
mem[11924] = 8'h02;
mem[11925] = 8'h95;
mem[11926] = 8'h0c;
mem[11927] = 8'ha9;
mem[11928] = 8'h00;
mem[11929] = 8'h48;
mem[11930] = 8'h28;
mem[11931] = 8'hd6;
mem[11932] = 8'h0c;
mem[11933] = 8'h08;
mem[11934] = 8'hb5;
mem[11935] = 8'h0c;
mem[11936] = 8'hdd;
mem[11937] = 8'h40;
mem[11938] = 8'h02;
mem[11939] = 8'hd0;
mem[11940] = 8'hfe;
mem[11941] = 8'h68;
mem[11942] = 8'h09;
mem[11943] = 8'h08;
mem[11944] = 8'h49;
mem[11945] = 8'h38;
mem[11946] = 8'hdd;
mem[11947] = 8'h45;
mem[11948] = 8'h02;
mem[11949] = 8'hd0;
mem[11950] = 8'hfe;
mem[11951] = 8'hb5;
mem[11952] = 8'h0c;
mem[11953] = 8'hca;
mem[11954] = 8'h30;
mem[11955] = 8'h08;
mem[11956] = 8'he0;
mem[11957] = 8'h01;
mem[11958] = 8'hd0;
mem[11959] = 8'hdd;
mem[11960] = 8'ha9;
mem[11961] = 8'h81;
mem[11962] = 8'hd0;
mem[11963] = 8'hd9;
mem[11964] = 8'ha2;
mem[11965] = 8'h00;
mem[11966] = 8'ha9;
mem[11967] = 8'h7e;
mem[11968] = 8'h95;
mem[11969] = 8'h0c;
mem[11970] = 8'ha9;
mem[11971] = 8'hff;
mem[11972] = 8'h48;
mem[11973] = 8'h28;
mem[11974] = 8'hf6;
mem[11975] = 8'h0c;
mem[11976] = 8'h08;
mem[11977] = 8'hb5;
mem[11978] = 8'h0c;
mem[11979] = 8'hdd;
mem[11980] = 8'h40;
mem[11981] = 8'h02;
mem[11982] = 8'hd0;
mem[11983] = 8'hfe;
mem[11984] = 8'h68;
mem[11985] = 8'h09;
mem[11986] = 8'h08;
mem[11987] = 8'h49;
mem[11988] = 8'h7d;
mem[11989] = 8'hdd;
mem[11990] = 8'h45;
mem[11991] = 8'h02;
mem[11992] = 8'hd0;
mem[11993] = 8'hfe;
mem[11994] = 8'hb5;
mem[11995] = 8'h0c;
mem[11996] = 8'he8;
mem[11997] = 8'he0;
mem[11998] = 8'h02;
mem[11999] = 8'hd0;
mem[12000] = 8'h02;
mem[12001] = 8'ha9;
mem[12002] = 8'hfe;
mem[12003] = 8'he0;
mem[12004] = 8'h05;
mem[12005] = 8'hd0;
mem[12006] = 8'hd9;
mem[12007] = 8'hca;
mem[12008] = 8'ha9;
mem[12009] = 8'h02;
mem[12010] = 8'h95;
mem[12011] = 8'h0c;
mem[12012] = 8'ha9;
mem[12013] = 8'hff;
mem[12014] = 8'h48;
mem[12015] = 8'h28;
mem[12016] = 8'hd6;
mem[12017] = 8'h0c;
mem[12018] = 8'h08;
mem[12019] = 8'hb5;
mem[12020] = 8'h0c;
mem[12021] = 8'hdd;
mem[12022] = 8'h40;
mem[12023] = 8'h02;
mem[12024] = 8'hd0;
mem[12025] = 8'hfe;
mem[12026] = 8'h68;
mem[12027] = 8'h09;
mem[12028] = 8'h08;
mem[12029] = 8'h49;
mem[12030] = 8'h7d;
mem[12031] = 8'hdd;
mem[12032] = 8'h45;
mem[12033] = 8'h02;
mem[12034] = 8'hd0;
mem[12035] = 8'hfe;
mem[12036] = 8'hb5;
mem[12037] = 8'h0c;
mem[12038] = 8'hca;
mem[12039] = 8'h30;
mem[12040] = 8'h08;
mem[12041] = 8'he0;
mem[12042] = 8'h01;
mem[12043] = 8'hd0;
mem[12044] = 8'hdd;
mem[12045] = 8'ha9;
mem[12046] = 8'h81;
mem[12047] = 8'hd0;
mem[12048] = 8'hd9;
mem[12049] = 8'had;
mem[12050] = 8'h00;
mem[12051] = 8'h02;
mem[12052] = 8'hc9;
mem[12053] = 8'h24;
mem[12054] = 8'hd0;
mem[12055] = 8'hfe;
mem[12056] = 8'ha9;
mem[12057] = 8'h25;
mem[12058] = 8'h8d;
mem[12059] = 8'h00;
mem[12060] = 8'h02;
mem[12061] = 8'ha2;
mem[12062] = 8'h00;
mem[12063] = 8'ha9;
mem[12064] = 8'h7e;
mem[12065] = 8'h9d;
mem[12066] = 8'h03;
mem[12067] = 8'h02;
mem[12068] = 8'ha9;
mem[12069] = 8'h00;
mem[12070] = 8'h48;
mem[12071] = 8'h28;
mem[12072] = 8'hfe;
mem[12073] = 8'h03;
mem[12074] = 8'h02;
mem[12075] = 8'h08;
mem[12076] = 8'hbd;
mem[12077] = 8'h03;
mem[12078] = 8'h02;
mem[12079] = 8'hdd;
mem[12080] = 8'h40;
mem[12081] = 8'h02;
mem[12082] = 8'hd0;
mem[12083] = 8'hfe;
mem[12084] = 8'h68;
mem[12085] = 8'h09;
mem[12086] = 8'h08;
mem[12087] = 8'h49;
mem[12088] = 8'h38;
mem[12089] = 8'hdd;
mem[12090] = 8'h45;
mem[12091] = 8'h02;
mem[12092] = 8'hd0;
mem[12093] = 8'hfe;
mem[12094] = 8'hbd;
mem[12095] = 8'h03;
mem[12096] = 8'h02;
mem[12097] = 8'he8;
mem[12098] = 8'he0;
mem[12099] = 8'h02;
mem[12100] = 8'hd0;
mem[12101] = 8'h02;
mem[12102] = 8'ha9;
mem[12103] = 8'hfe;
mem[12104] = 8'he0;
mem[12105] = 8'h05;
mem[12106] = 8'hd0;
mem[12107] = 8'hd5;
mem[12108] = 8'hca;
mem[12109] = 8'ha9;
mem[12110] = 8'h02;
mem[12111] = 8'h9d;
mem[12112] = 8'h03;
mem[12113] = 8'h02;
mem[12114] = 8'ha9;
mem[12115] = 8'h00;
mem[12116] = 8'h48;
mem[12117] = 8'h28;
mem[12118] = 8'hde;
mem[12119] = 8'h03;
mem[12120] = 8'h02;
mem[12121] = 8'h08;
mem[12122] = 8'hbd;
mem[12123] = 8'h03;
mem[12124] = 8'h02;
mem[12125] = 8'hdd;
mem[12126] = 8'h40;
mem[12127] = 8'h02;
mem[12128] = 8'hd0;
mem[12129] = 8'hfe;
mem[12130] = 8'h68;
mem[12131] = 8'h09;
mem[12132] = 8'h08;
mem[12133] = 8'h49;
mem[12134] = 8'h38;
mem[12135] = 8'hdd;
mem[12136] = 8'h45;
mem[12137] = 8'h02;
mem[12138] = 8'hd0;
mem[12139] = 8'hfe;
mem[12140] = 8'hbd;
mem[12141] = 8'h03;
mem[12142] = 8'h02;
mem[12143] = 8'hca;
mem[12144] = 8'h30;
mem[12145] = 8'h08;
mem[12146] = 8'he0;
mem[12147] = 8'h01;
mem[12148] = 8'hd0;
mem[12149] = 8'hd9;
mem[12150] = 8'ha9;
mem[12151] = 8'h81;
mem[12152] = 8'hd0;
mem[12153] = 8'hd5;
mem[12154] = 8'ha2;
mem[12155] = 8'h00;
mem[12156] = 8'ha9;
mem[12157] = 8'h7e;
mem[12158] = 8'h9d;
mem[12159] = 8'h03;
mem[12160] = 8'h02;
mem[12161] = 8'ha9;
mem[12162] = 8'hff;
mem[12163] = 8'h48;
mem[12164] = 8'h28;
mem[12165] = 8'hfe;
mem[12166] = 8'h03;
mem[12167] = 8'h02;
mem[12168] = 8'h08;
mem[12169] = 8'hbd;
mem[12170] = 8'h03;
mem[12171] = 8'h02;
mem[12172] = 8'hdd;
mem[12173] = 8'h40;
mem[12174] = 8'h02;
mem[12175] = 8'hd0;
mem[12176] = 8'hfe;
mem[12177] = 8'h68;
mem[12178] = 8'h09;
mem[12179] = 8'h08;
mem[12180] = 8'h49;
mem[12181] = 8'h7d;
mem[12182] = 8'hdd;
mem[12183] = 8'h45;
mem[12184] = 8'h02;
mem[12185] = 8'hd0;
mem[12186] = 8'hfe;
mem[12187] = 8'hbd;
mem[12188] = 8'h03;
mem[12189] = 8'h02;
mem[12190] = 8'he8;
mem[12191] = 8'he0;
mem[12192] = 8'h02;
mem[12193] = 8'hd0;
mem[12194] = 8'h02;
mem[12195] = 8'ha9;
mem[12196] = 8'hfe;
mem[12197] = 8'he0;
mem[12198] = 8'h05;
mem[12199] = 8'hd0;
mem[12200] = 8'hd5;
mem[12201] = 8'hca;
mem[12202] = 8'ha9;
mem[12203] = 8'h02;
mem[12204] = 8'h9d;
mem[12205] = 8'h03;
mem[12206] = 8'h02;
mem[12207] = 8'ha9;
mem[12208] = 8'hff;
mem[12209] = 8'h48;
mem[12210] = 8'h28;
mem[12211] = 8'hde;
mem[12212] = 8'h03;
mem[12213] = 8'h02;
mem[12214] = 8'h08;
mem[12215] = 8'hbd;
mem[12216] = 8'h03;
mem[12217] = 8'h02;
mem[12218] = 8'hdd;
mem[12219] = 8'h40;
mem[12220] = 8'h02;
mem[12221] = 8'hd0;
mem[12222] = 8'hfe;
mem[12223] = 8'h68;
mem[12224] = 8'h09;
mem[12225] = 8'h08;
mem[12226] = 8'h49;
mem[12227] = 8'h7d;
mem[12228] = 8'hdd;
mem[12229] = 8'h45;
mem[12230] = 8'h02;
mem[12231] = 8'hd0;
mem[12232] = 8'hfe;
mem[12233] = 8'hbd;
mem[12234] = 8'h03;
mem[12235] = 8'h02;
mem[12236] = 8'hca;
mem[12237] = 8'h30;
mem[12238] = 8'h08;
mem[12239] = 8'he0;
mem[12240] = 8'h01;
mem[12241] = 8'hd0;
mem[12242] = 8'hd9;
mem[12243] = 8'ha9;
mem[12244] = 8'h81;
mem[12245] = 8'hd0;
mem[12246] = 8'hd5;
mem[12247] = 8'had;
mem[12248] = 8'h00;
mem[12249] = 8'h02;
mem[12250] = 8'hc9;
mem[12251] = 8'h25;
mem[12252] = 8'hd0;
mem[12253] = 8'hfe;
mem[12254] = 8'ha9;
mem[12255] = 8'h26;
mem[12256] = 8'h8d;
mem[12257] = 8'h00;
mem[12258] = 8'h02;
mem[12259] = 8'ha2;
mem[12260] = 8'h03;
mem[12261] = 8'hb5;
mem[12262] = 8'h1c;
mem[12263] = 8'h8d;
mem[12264] = 8'h09;
mem[12265] = 8'h02;
mem[12266] = 8'ha9;
mem[12267] = 8'h00;
mem[12268] = 8'h48;
mem[12269] = 8'hbd;
mem[12270] = 8'h5a;
mem[12271] = 8'h02;
mem[12272] = 8'h28;
mem[12273] = 8'h20;
mem[12274] = 8'h08;
mem[12275] = 8'h02;
mem[12276] = 8'h08;
mem[12277] = 8'hdd;
mem[12278] = 8'h62;
mem[12279] = 8'h02;
mem[12280] = 8'hd0;
mem[12281] = 8'hfe;
mem[12282] = 8'h68;
mem[12283] = 8'h09;
mem[12284] = 8'h08;
mem[12285] = 8'h49;
mem[12286] = 8'h38;
mem[12287] = 8'hdd;
mem[12288] = 8'h66;
mem[12289] = 8'h02;
mem[12290] = 8'hd0;
mem[12291] = 8'hfe;
mem[12292] = 8'hca;
mem[12293] = 8'h10;
mem[12294] = 8'hde;
mem[12295] = 8'ha2;
mem[12296] = 8'h03;
mem[12297] = 8'hb5;
mem[12298] = 8'h1c;
mem[12299] = 8'h8d;
mem[12300] = 8'h09;
mem[12301] = 8'h02;
mem[12302] = 8'ha9;
mem[12303] = 8'hff;
mem[12304] = 8'h48;
mem[12305] = 8'hbd;
mem[12306] = 8'h5a;
mem[12307] = 8'h02;
mem[12308] = 8'h28;
mem[12309] = 8'h20;
mem[12310] = 8'h08;
mem[12311] = 8'h02;
mem[12312] = 8'h08;
mem[12313] = 8'hdd;
mem[12314] = 8'h62;
mem[12315] = 8'h02;
mem[12316] = 8'hd0;
mem[12317] = 8'hfe;
mem[12318] = 8'h68;
mem[12319] = 8'h09;
mem[12320] = 8'h08;
mem[12321] = 8'h49;
mem[12322] = 8'h7d;
mem[12323] = 8'hdd;
mem[12324] = 8'h66;
mem[12325] = 8'h02;
mem[12326] = 8'hd0;
mem[12327] = 8'hfe;
mem[12328] = 8'hca;
mem[12329] = 8'h10;
mem[12330] = 8'hde;
mem[12331] = 8'ha2;
mem[12332] = 8'h03;
mem[12333] = 8'hb5;
mem[12334] = 8'h1c;
mem[12335] = 8'h85;
mem[12336] = 8'h0c;
mem[12337] = 8'ha9;
mem[12338] = 8'h00;
mem[12339] = 8'h48;
mem[12340] = 8'hbd;
mem[12341] = 8'h5a;
mem[12342] = 8'h02;
mem[12343] = 8'h28;
mem[12344] = 8'h25;
mem[12345] = 8'h0c;
mem[12346] = 8'h08;
mem[12347] = 8'hdd;
mem[12348] = 8'h62;
mem[12349] = 8'h02;
mem[12350] = 8'hd0;
mem[12351] = 8'hfe;
mem[12352] = 8'h68;
mem[12353] = 8'h09;
mem[12354] = 8'h08;
mem[12355] = 8'h49;
mem[12356] = 8'h38;
mem[12357] = 8'hdd;
mem[12358] = 8'h66;
mem[12359] = 8'h02;
mem[12360] = 8'hd0;
mem[12361] = 8'hfe;
mem[12362] = 8'hca;
mem[12363] = 8'h10;
mem[12364] = 8'he0;
mem[12365] = 8'ha2;
mem[12366] = 8'h03;
mem[12367] = 8'hb5;
mem[12368] = 8'h1c;
mem[12369] = 8'h85;
mem[12370] = 8'h0c;
mem[12371] = 8'ha9;
mem[12372] = 8'hff;
mem[12373] = 8'h48;
mem[12374] = 8'hbd;
mem[12375] = 8'h5a;
mem[12376] = 8'h02;
mem[12377] = 8'h28;
mem[12378] = 8'h25;
mem[12379] = 8'h0c;
mem[12380] = 8'h08;
mem[12381] = 8'hdd;
mem[12382] = 8'h62;
mem[12383] = 8'h02;
mem[12384] = 8'hd0;
mem[12385] = 8'hfe;
mem[12386] = 8'h68;
mem[12387] = 8'h09;
mem[12388] = 8'h08;
mem[12389] = 8'h49;
mem[12390] = 8'h7d;
mem[12391] = 8'hdd;
mem[12392] = 8'h66;
mem[12393] = 8'h02;
mem[12394] = 8'hd0;
mem[12395] = 8'hfe;
mem[12396] = 8'hca;
mem[12397] = 8'h10;
mem[12398] = 8'he0;
mem[12399] = 8'ha2;
mem[12400] = 8'h03;
mem[12401] = 8'hb5;
mem[12402] = 8'h1c;
mem[12403] = 8'h8d;
mem[12404] = 8'h03;
mem[12405] = 8'h02;
mem[12406] = 8'ha9;
mem[12407] = 8'h00;
mem[12408] = 8'h48;
mem[12409] = 8'hbd;
mem[12410] = 8'h5a;
mem[12411] = 8'h02;
mem[12412] = 8'h28;
mem[12413] = 8'h2d;
mem[12414] = 8'h03;
mem[12415] = 8'h02;
mem[12416] = 8'h08;
mem[12417] = 8'hdd;
mem[12418] = 8'h62;
mem[12419] = 8'h02;
mem[12420] = 8'hd0;
mem[12421] = 8'hfe;
mem[12422] = 8'h68;
mem[12423] = 8'h09;
mem[12424] = 8'h08;
mem[12425] = 8'h49;
mem[12426] = 8'h38;
mem[12427] = 8'hdd;
mem[12428] = 8'h66;
mem[12429] = 8'h02;
mem[12430] = 8'hd0;
mem[12431] = 8'hfe;
mem[12432] = 8'hca;
mem[12433] = 8'h10;
mem[12434] = 8'hde;
mem[12435] = 8'ha2;
mem[12436] = 8'h03;
mem[12437] = 8'hb5;
mem[12438] = 8'h1c;
mem[12439] = 8'h8d;
mem[12440] = 8'h03;
mem[12441] = 8'h02;
mem[12442] = 8'ha9;
mem[12443] = 8'hff;
mem[12444] = 8'h48;
mem[12445] = 8'hbd;
mem[12446] = 8'h5a;
mem[12447] = 8'h02;
mem[12448] = 8'h28;
mem[12449] = 8'h2d;
mem[12450] = 8'h03;
mem[12451] = 8'h02;
mem[12452] = 8'h08;
mem[12453] = 8'hdd;
mem[12454] = 8'h62;
mem[12455] = 8'h02;
mem[12456] = 8'hd0;
mem[12457] = 8'hfe;
mem[12458] = 8'h68;
mem[12459] = 8'h09;
mem[12460] = 8'h08;
mem[12461] = 8'h49;
mem[12462] = 8'h7d;
mem[12463] = 8'hdd;
mem[12464] = 8'h66;
mem[12465] = 8'h02;
mem[12466] = 8'hd0;
mem[12467] = 8'hfe;
mem[12468] = 8'hca;
mem[12469] = 8'h10;
mem[12470] = 8'h02;
mem[12471] = 8'ha2;
mem[12472] = 8'h03;
mem[12473] = 8'ha9;
mem[12474] = 8'h00;
mem[12475] = 8'h48;
mem[12476] = 8'hbd;
mem[12477] = 8'h5a;
mem[12478] = 8'h02;
mem[12479] = 8'h28;
mem[12480] = 8'h35;
mem[12481] = 8'h1c;
mem[12482] = 8'h08;
mem[12483] = 8'hdd;
mem[12484] = 8'h62;
mem[12485] = 8'h02;
mem[12486] = 8'hd0;
mem[12487] = 8'hfe;
mem[12488] = 8'h68;
mem[12489] = 8'h09;
mem[12490] = 8'h08;
mem[12491] = 8'h49;
mem[12492] = 8'h38;
mem[12493] = 8'hdd;
mem[12494] = 8'h66;
mem[12495] = 8'h02;
mem[12496] = 8'hd0;
mem[12497] = 8'hfe;
mem[12498] = 8'hca;
mem[12499] = 8'h10;
mem[12500] = 8'he4;
mem[12501] = 8'ha2;
mem[12502] = 8'h03;
mem[12503] = 8'ha9;
mem[12504] = 8'hff;
mem[12505] = 8'h48;
mem[12506] = 8'hbd;
mem[12507] = 8'h5a;
mem[12508] = 8'h02;
mem[12509] = 8'h28;
mem[12510] = 8'h35;
mem[12511] = 8'h1c;
mem[12512] = 8'h08;
mem[12513] = 8'hdd;
mem[12514] = 8'h62;
mem[12515] = 8'h02;
mem[12516] = 8'hd0;
mem[12517] = 8'hfe;
mem[12518] = 8'h68;
mem[12519] = 8'h09;
mem[12520] = 8'h08;
mem[12521] = 8'h49;
mem[12522] = 8'h7d;
mem[12523] = 8'hdd;
mem[12524] = 8'h66;
mem[12525] = 8'h02;
mem[12526] = 8'hd0;
mem[12527] = 8'hfe;
mem[12528] = 8'hca;
mem[12529] = 8'h10;
mem[12530] = 8'he4;
mem[12531] = 8'ha2;
mem[12532] = 8'h03;
mem[12533] = 8'ha9;
mem[12534] = 8'h00;
mem[12535] = 8'h48;
mem[12536] = 8'hbd;
mem[12537] = 8'h5a;
mem[12538] = 8'h02;
mem[12539] = 8'h28;
mem[12540] = 8'h3d;
mem[12541] = 8'h4e;
mem[12542] = 8'h02;
mem[12543] = 8'h08;
mem[12544] = 8'hdd;
mem[12545] = 8'h62;
mem[12546] = 8'h02;
mem[12547] = 8'hd0;
mem[12548] = 8'hfe;
mem[12549] = 8'h68;
mem[12550] = 8'h09;
mem[12551] = 8'h08;
mem[12552] = 8'h49;
mem[12553] = 8'h38;
mem[12554] = 8'hdd;
mem[12555] = 8'h66;
mem[12556] = 8'h02;
mem[12557] = 8'hd0;
mem[12558] = 8'hfe;
mem[12559] = 8'hca;
mem[12560] = 8'h10;
mem[12561] = 8'he3;
mem[12562] = 8'ha2;
mem[12563] = 8'h03;
mem[12564] = 8'ha9;
mem[12565] = 8'hff;
mem[12566] = 8'h48;
mem[12567] = 8'hbd;
mem[12568] = 8'h5a;
mem[12569] = 8'h02;
mem[12570] = 8'h28;
mem[12571] = 8'h3d;
mem[12572] = 8'h4e;
mem[12573] = 8'h02;
mem[12574] = 8'h08;
mem[12575] = 8'hdd;
mem[12576] = 8'h62;
mem[12577] = 8'h02;
mem[12578] = 8'hd0;
mem[12579] = 8'hfe;
mem[12580] = 8'h68;
mem[12581] = 8'h09;
mem[12582] = 8'h08;
mem[12583] = 8'h49;
mem[12584] = 8'h7d;
mem[12585] = 8'hdd;
mem[12586] = 8'h66;
mem[12587] = 8'h02;
mem[12588] = 8'hd0;
mem[12589] = 8'hfe;
mem[12590] = 8'hca;
mem[12591] = 8'h10;
mem[12592] = 8'he3;
mem[12593] = 8'ha0;
mem[12594] = 8'h03;
mem[12595] = 8'ha9;
mem[12596] = 8'h00;
mem[12597] = 8'h48;
mem[12598] = 8'hb9;
mem[12599] = 8'h5a;
mem[12600] = 8'h02;
mem[12601] = 8'h28;
mem[12602] = 8'h39;
mem[12603] = 8'h4e;
mem[12604] = 8'h02;
mem[12605] = 8'h08;
mem[12606] = 8'hd9;
mem[12607] = 8'h62;
mem[12608] = 8'h02;
mem[12609] = 8'hd0;
mem[12610] = 8'hfe;
mem[12611] = 8'h68;
mem[12612] = 8'h09;
mem[12613] = 8'h08;
mem[12614] = 8'h49;
mem[12615] = 8'h38;
mem[12616] = 8'hd9;
mem[12617] = 8'h66;
mem[12618] = 8'h02;
mem[12619] = 8'hd0;
mem[12620] = 8'hfe;
mem[12621] = 8'h88;
mem[12622] = 8'h10;
mem[12623] = 8'he3;
mem[12624] = 8'ha0;
mem[12625] = 8'h03;
mem[12626] = 8'ha9;
mem[12627] = 8'hff;
mem[12628] = 8'h48;
mem[12629] = 8'hb9;
mem[12630] = 8'h5a;
mem[12631] = 8'h02;
mem[12632] = 8'h28;
mem[12633] = 8'h39;
mem[12634] = 8'h4e;
mem[12635] = 8'h02;
mem[12636] = 8'h08;
mem[12637] = 8'hd9;
mem[12638] = 8'h62;
mem[12639] = 8'h02;
mem[12640] = 8'hd0;
mem[12641] = 8'hfe;
mem[12642] = 8'h68;
mem[12643] = 8'h09;
mem[12644] = 8'h08;
mem[12645] = 8'h49;
mem[12646] = 8'h7d;
mem[12647] = 8'hd9;
mem[12648] = 8'h66;
mem[12649] = 8'h02;
mem[12650] = 8'hd0;
mem[12651] = 8'hfe;
mem[12652] = 8'h88;
mem[12653] = 8'h10;
mem[12654] = 8'he3;
mem[12655] = 8'ha2;
mem[12656] = 8'h06;
mem[12657] = 8'ha0;
mem[12658] = 8'h03;
mem[12659] = 8'ha9;
mem[12660] = 8'h00;
mem[12661] = 8'h48;
mem[12662] = 8'hb9;
mem[12663] = 8'h5a;
mem[12664] = 8'h02;
mem[12665] = 8'h28;
mem[12666] = 8'h21;
mem[12667] = 8'h3a;
mem[12668] = 8'h08;
mem[12669] = 8'hd9;
mem[12670] = 8'h62;
mem[12671] = 8'h02;
mem[12672] = 8'hd0;
mem[12673] = 8'hfe;
mem[12674] = 8'h68;
mem[12675] = 8'h09;
mem[12676] = 8'h08;
mem[12677] = 8'h49;
mem[12678] = 8'h38;
mem[12679] = 8'hd9;
mem[12680] = 8'h66;
mem[12681] = 8'h02;
mem[12682] = 8'hd0;
mem[12683] = 8'hfe;
mem[12684] = 8'hca;
mem[12685] = 8'hca;
mem[12686] = 8'h88;
mem[12687] = 8'h10;
mem[12688] = 8'he2;
mem[12689] = 8'ha2;
mem[12690] = 8'h06;
mem[12691] = 8'ha0;
mem[12692] = 8'h03;
mem[12693] = 8'ha9;
mem[12694] = 8'hff;
mem[12695] = 8'h48;
mem[12696] = 8'hb9;
mem[12697] = 8'h5a;
mem[12698] = 8'h02;
mem[12699] = 8'h28;
mem[12700] = 8'h21;
mem[12701] = 8'h3a;
mem[12702] = 8'h08;
mem[12703] = 8'hd9;
mem[12704] = 8'h62;
mem[12705] = 8'h02;
mem[12706] = 8'hd0;
mem[12707] = 8'hfe;
mem[12708] = 8'h68;
mem[12709] = 8'h09;
mem[12710] = 8'h08;
mem[12711] = 8'h49;
mem[12712] = 8'h7d;
mem[12713] = 8'hd9;
mem[12714] = 8'h66;
mem[12715] = 8'h02;
mem[12716] = 8'hd0;
mem[12717] = 8'hfe;
mem[12718] = 8'hca;
mem[12719] = 8'hca;
mem[12720] = 8'h88;
mem[12721] = 8'h10;
mem[12722] = 8'he2;
mem[12723] = 8'ha0;
mem[12724] = 8'h03;
mem[12725] = 8'ha9;
mem[12726] = 8'h00;
mem[12727] = 8'h48;
mem[12728] = 8'hb9;
mem[12729] = 8'h5a;
mem[12730] = 8'h02;
mem[12731] = 8'h28;
mem[12732] = 8'h31;
mem[12733] = 8'h3a;
mem[12734] = 8'h08;
mem[12735] = 8'hd9;
mem[12736] = 8'h62;
mem[12737] = 8'h02;
mem[12738] = 8'hd0;
mem[12739] = 8'hfe;
mem[12740] = 8'h68;
mem[12741] = 8'h09;
mem[12742] = 8'h08;
mem[12743] = 8'h49;
mem[12744] = 8'h38;
mem[12745] = 8'hd9;
mem[12746] = 8'h66;
mem[12747] = 8'h02;
mem[12748] = 8'hd0;
mem[12749] = 8'hfe;
mem[12750] = 8'h88;
mem[12751] = 8'h10;
mem[12752] = 8'he4;
mem[12753] = 8'ha0;
mem[12754] = 8'h03;
mem[12755] = 8'ha9;
mem[12756] = 8'hff;
mem[12757] = 8'h48;
mem[12758] = 8'hb9;
mem[12759] = 8'h5a;
mem[12760] = 8'h02;
mem[12761] = 8'h28;
mem[12762] = 8'h31;
mem[12763] = 8'h3a;
mem[12764] = 8'h08;
mem[12765] = 8'hd9;
mem[12766] = 8'h62;
mem[12767] = 8'h02;
mem[12768] = 8'hd0;
mem[12769] = 8'hfe;
mem[12770] = 8'h68;
mem[12771] = 8'h09;
mem[12772] = 8'h08;
mem[12773] = 8'h49;
mem[12774] = 8'h7d;
mem[12775] = 8'hd9;
mem[12776] = 8'h66;
mem[12777] = 8'h02;
mem[12778] = 8'hd0;
mem[12779] = 8'hfe;
mem[12780] = 8'h88;
mem[12781] = 8'h10;
mem[12782] = 8'he4;
mem[12783] = 8'had;
mem[12784] = 8'h00;
mem[12785] = 8'h02;
mem[12786] = 8'hc9;
mem[12787] = 8'h26;
mem[12788] = 8'hd0;
mem[12789] = 8'hfe;
mem[12790] = 8'ha9;
mem[12791] = 8'h27;
mem[12792] = 8'h8d;
mem[12793] = 8'h00;
mem[12794] = 8'h02;
mem[12795] = 8'ha2;
mem[12796] = 8'h03;
mem[12797] = 8'hb5;
mem[12798] = 8'h20;
mem[12799] = 8'h8d;
mem[12800] = 8'h0c;
mem[12801] = 8'h02;
mem[12802] = 8'ha9;
mem[12803] = 8'h00;
mem[12804] = 8'h48;
mem[12805] = 8'hbd;
mem[12806] = 8'h5e;
mem[12807] = 8'h02;
mem[12808] = 8'h28;
mem[12809] = 8'h20;
mem[12810] = 8'h0b;
mem[12811] = 8'h02;
mem[12812] = 8'h08;
mem[12813] = 8'hdd;
mem[12814] = 8'h62;
mem[12815] = 8'h02;
mem[12816] = 8'hd0;
mem[12817] = 8'hfe;
mem[12818] = 8'h68;
mem[12819] = 8'h09;
mem[12820] = 8'h08;
mem[12821] = 8'h49;
mem[12822] = 8'h38;
mem[12823] = 8'hdd;
mem[12824] = 8'h66;
mem[12825] = 8'h02;
mem[12826] = 8'hd0;
mem[12827] = 8'hfe;
mem[12828] = 8'hca;
mem[12829] = 8'h10;
mem[12830] = 8'hde;
mem[12831] = 8'ha2;
mem[12832] = 8'h03;
mem[12833] = 8'hb5;
mem[12834] = 8'h20;
mem[12835] = 8'h8d;
mem[12836] = 8'h0c;
mem[12837] = 8'h02;
mem[12838] = 8'ha9;
mem[12839] = 8'hff;
mem[12840] = 8'h48;
mem[12841] = 8'hbd;
mem[12842] = 8'h5e;
mem[12843] = 8'h02;
mem[12844] = 8'h28;
mem[12845] = 8'h20;
mem[12846] = 8'h0b;
mem[12847] = 8'h02;
mem[12848] = 8'h08;
mem[12849] = 8'hdd;
mem[12850] = 8'h62;
mem[12851] = 8'h02;
mem[12852] = 8'hd0;
mem[12853] = 8'hfe;
mem[12854] = 8'h68;
mem[12855] = 8'h09;
mem[12856] = 8'h08;
mem[12857] = 8'h49;
mem[12858] = 8'h7d;
mem[12859] = 8'hdd;
mem[12860] = 8'h66;
mem[12861] = 8'h02;
mem[12862] = 8'hd0;
mem[12863] = 8'hfe;
mem[12864] = 8'hca;
mem[12865] = 8'h10;
mem[12866] = 8'hde;
mem[12867] = 8'ha2;
mem[12868] = 8'h03;
mem[12869] = 8'hb5;
mem[12870] = 8'h20;
mem[12871] = 8'h85;
mem[12872] = 8'h0c;
mem[12873] = 8'ha9;
mem[12874] = 8'h00;
mem[12875] = 8'h48;
mem[12876] = 8'hbd;
mem[12877] = 8'h5e;
mem[12878] = 8'h02;
mem[12879] = 8'h28;
mem[12880] = 8'h45;
mem[12881] = 8'h0c;
mem[12882] = 8'h08;
mem[12883] = 8'hdd;
mem[12884] = 8'h62;
mem[12885] = 8'h02;
mem[12886] = 8'hd0;
mem[12887] = 8'hfe;
mem[12888] = 8'h68;
mem[12889] = 8'h09;
mem[12890] = 8'h08;
mem[12891] = 8'h49;
mem[12892] = 8'h38;
mem[12893] = 8'hdd;
mem[12894] = 8'h66;
mem[12895] = 8'h02;
mem[12896] = 8'hd0;
mem[12897] = 8'hfe;
mem[12898] = 8'hca;
mem[12899] = 8'h10;
mem[12900] = 8'he0;
mem[12901] = 8'ha2;
mem[12902] = 8'h03;
mem[12903] = 8'hb5;
mem[12904] = 8'h20;
mem[12905] = 8'h85;
mem[12906] = 8'h0c;
mem[12907] = 8'ha9;
mem[12908] = 8'hff;
mem[12909] = 8'h48;
mem[12910] = 8'hbd;
mem[12911] = 8'h5e;
mem[12912] = 8'h02;
mem[12913] = 8'h28;
mem[12914] = 8'h45;
mem[12915] = 8'h0c;
mem[12916] = 8'h08;
mem[12917] = 8'hdd;
mem[12918] = 8'h62;
mem[12919] = 8'h02;
mem[12920] = 8'hd0;
mem[12921] = 8'hfe;
mem[12922] = 8'h68;
mem[12923] = 8'h09;
mem[12924] = 8'h08;
mem[12925] = 8'h49;
mem[12926] = 8'h7d;
mem[12927] = 8'hdd;
mem[12928] = 8'h66;
mem[12929] = 8'h02;
mem[12930] = 8'hd0;
mem[12931] = 8'hfe;
mem[12932] = 8'hca;
mem[12933] = 8'h10;
mem[12934] = 8'he0;
mem[12935] = 8'ha2;
mem[12936] = 8'h03;
mem[12937] = 8'hb5;
mem[12938] = 8'h20;
mem[12939] = 8'h8d;
mem[12940] = 8'h03;
mem[12941] = 8'h02;
mem[12942] = 8'ha9;
mem[12943] = 8'h00;
mem[12944] = 8'h48;
mem[12945] = 8'hbd;
mem[12946] = 8'h5e;
mem[12947] = 8'h02;
mem[12948] = 8'h28;
mem[12949] = 8'h4d;
mem[12950] = 8'h03;
mem[12951] = 8'h02;
mem[12952] = 8'h08;
mem[12953] = 8'hdd;
mem[12954] = 8'h62;
mem[12955] = 8'h02;
mem[12956] = 8'hd0;
mem[12957] = 8'hfe;
mem[12958] = 8'h68;
mem[12959] = 8'h09;
mem[12960] = 8'h08;
mem[12961] = 8'h49;
mem[12962] = 8'h38;
mem[12963] = 8'hdd;
mem[12964] = 8'h66;
mem[12965] = 8'h02;
mem[12966] = 8'hd0;
mem[12967] = 8'hfe;
mem[12968] = 8'hca;
mem[12969] = 8'h10;
mem[12970] = 8'hde;
mem[12971] = 8'ha2;
mem[12972] = 8'h03;
mem[12973] = 8'hb5;
mem[12974] = 8'h20;
mem[12975] = 8'h8d;
mem[12976] = 8'h03;
mem[12977] = 8'h02;
mem[12978] = 8'ha9;
mem[12979] = 8'hff;
mem[12980] = 8'h48;
mem[12981] = 8'hbd;
mem[12982] = 8'h5e;
mem[12983] = 8'h02;
mem[12984] = 8'h28;
mem[12985] = 8'h4d;
mem[12986] = 8'h03;
mem[12987] = 8'h02;
mem[12988] = 8'h08;
mem[12989] = 8'hdd;
mem[12990] = 8'h62;
mem[12991] = 8'h02;
mem[12992] = 8'hd0;
mem[12993] = 8'hfe;
mem[12994] = 8'h68;
mem[12995] = 8'h09;
mem[12996] = 8'h08;
mem[12997] = 8'h49;
mem[12998] = 8'h7d;
mem[12999] = 8'hdd;
mem[13000] = 8'h66;
mem[13001] = 8'h02;
mem[13002] = 8'hd0;
mem[13003] = 8'hfe;
mem[13004] = 8'hca;
mem[13005] = 8'h10;
mem[13006] = 8'h02;
mem[13007] = 8'ha2;
mem[13008] = 8'h03;
mem[13009] = 8'ha9;
mem[13010] = 8'h00;
mem[13011] = 8'h48;
mem[13012] = 8'hbd;
mem[13013] = 8'h5e;
mem[13014] = 8'h02;
mem[13015] = 8'h28;
mem[13016] = 8'h55;
mem[13017] = 8'h20;
mem[13018] = 8'h08;
mem[13019] = 8'hdd;
mem[13020] = 8'h62;
mem[13021] = 8'h02;
mem[13022] = 8'hd0;
mem[13023] = 8'hfe;
mem[13024] = 8'h68;
mem[13025] = 8'h09;
mem[13026] = 8'h08;
mem[13027] = 8'h49;
mem[13028] = 8'h38;
mem[13029] = 8'hdd;
mem[13030] = 8'h66;
mem[13031] = 8'h02;
mem[13032] = 8'hd0;
mem[13033] = 8'hfe;
mem[13034] = 8'hca;
mem[13035] = 8'h10;
mem[13036] = 8'he4;
mem[13037] = 8'ha2;
mem[13038] = 8'h03;
mem[13039] = 8'ha9;
mem[13040] = 8'hff;
mem[13041] = 8'h48;
mem[13042] = 8'hbd;
mem[13043] = 8'h5e;
mem[13044] = 8'h02;
mem[13045] = 8'h28;
mem[13046] = 8'h55;
mem[13047] = 8'h20;
mem[13048] = 8'h08;
mem[13049] = 8'hdd;
mem[13050] = 8'h62;
mem[13051] = 8'h02;
mem[13052] = 8'hd0;
mem[13053] = 8'hfe;
mem[13054] = 8'h68;
mem[13055] = 8'h09;
mem[13056] = 8'h08;
mem[13057] = 8'h49;
mem[13058] = 8'h7d;
mem[13059] = 8'hdd;
mem[13060] = 8'h66;
mem[13061] = 8'h02;
mem[13062] = 8'hd0;
mem[13063] = 8'hfe;
mem[13064] = 8'hca;
mem[13065] = 8'h10;
mem[13066] = 8'he4;
mem[13067] = 8'ha2;
mem[13068] = 8'h03;
mem[13069] = 8'ha9;
mem[13070] = 8'h00;
mem[13071] = 8'h48;
mem[13072] = 8'hbd;
mem[13073] = 8'h5e;
mem[13074] = 8'h02;
mem[13075] = 8'h28;
mem[13076] = 8'h5d;
mem[13077] = 8'h52;
mem[13078] = 8'h02;
mem[13079] = 8'h08;
mem[13080] = 8'hdd;
mem[13081] = 8'h62;
mem[13082] = 8'h02;
mem[13083] = 8'hd0;
mem[13084] = 8'hfe;
mem[13085] = 8'h68;
mem[13086] = 8'h09;
mem[13087] = 8'h08;
mem[13088] = 8'h49;
mem[13089] = 8'h38;
mem[13090] = 8'hdd;
mem[13091] = 8'h66;
mem[13092] = 8'h02;
mem[13093] = 8'hd0;
mem[13094] = 8'hfe;
mem[13095] = 8'hca;
mem[13096] = 8'h10;
mem[13097] = 8'he3;
mem[13098] = 8'ha2;
mem[13099] = 8'h03;
mem[13100] = 8'ha9;
mem[13101] = 8'hff;
mem[13102] = 8'h48;
mem[13103] = 8'hbd;
mem[13104] = 8'h5e;
mem[13105] = 8'h02;
mem[13106] = 8'h28;
mem[13107] = 8'h5d;
mem[13108] = 8'h52;
mem[13109] = 8'h02;
mem[13110] = 8'h08;
mem[13111] = 8'hdd;
mem[13112] = 8'h62;
mem[13113] = 8'h02;
mem[13114] = 8'hd0;
mem[13115] = 8'hfe;
mem[13116] = 8'h68;
mem[13117] = 8'h09;
mem[13118] = 8'h08;
mem[13119] = 8'h49;
mem[13120] = 8'h7d;
mem[13121] = 8'hdd;
mem[13122] = 8'h66;
mem[13123] = 8'h02;
mem[13124] = 8'hd0;
mem[13125] = 8'hfe;
mem[13126] = 8'hca;
mem[13127] = 8'h10;
mem[13128] = 8'he3;
mem[13129] = 8'ha0;
mem[13130] = 8'h03;
mem[13131] = 8'ha9;
mem[13132] = 8'h00;
mem[13133] = 8'h48;
mem[13134] = 8'hb9;
mem[13135] = 8'h5e;
mem[13136] = 8'h02;
mem[13137] = 8'h28;
mem[13138] = 8'h59;
mem[13139] = 8'h52;
mem[13140] = 8'h02;
mem[13141] = 8'h08;
mem[13142] = 8'hd9;
mem[13143] = 8'h62;
mem[13144] = 8'h02;
mem[13145] = 8'hd0;
mem[13146] = 8'hfe;
mem[13147] = 8'h68;
mem[13148] = 8'h09;
mem[13149] = 8'h08;
mem[13150] = 8'h49;
mem[13151] = 8'h38;
mem[13152] = 8'hd9;
mem[13153] = 8'h66;
mem[13154] = 8'h02;
mem[13155] = 8'hd0;
mem[13156] = 8'hfe;
mem[13157] = 8'h88;
mem[13158] = 8'h10;
mem[13159] = 8'he3;
mem[13160] = 8'ha0;
mem[13161] = 8'h03;
mem[13162] = 8'ha9;
mem[13163] = 8'hff;
mem[13164] = 8'h48;
mem[13165] = 8'hb9;
mem[13166] = 8'h5e;
mem[13167] = 8'h02;
mem[13168] = 8'h28;
mem[13169] = 8'h59;
mem[13170] = 8'h52;
mem[13171] = 8'h02;
mem[13172] = 8'h08;
mem[13173] = 8'hd9;
mem[13174] = 8'h62;
mem[13175] = 8'h02;
mem[13176] = 8'hd0;
mem[13177] = 8'hfe;
mem[13178] = 8'h68;
mem[13179] = 8'h09;
mem[13180] = 8'h08;
mem[13181] = 8'h49;
mem[13182] = 8'h7d;
mem[13183] = 8'hd9;
mem[13184] = 8'h66;
mem[13185] = 8'h02;
mem[13186] = 8'hd0;
mem[13187] = 8'hfe;
mem[13188] = 8'h88;
mem[13189] = 8'h10;
mem[13190] = 8'he3;
mem[13191] = 8'ha2;
mem[13192] = 8'h06;
mem[13193] = 8'ha0;
mem[13194] = 8'h03;
mem[13195] = 8'ha9;
mem[13196] = 8'h00;
mem[13197] = 8'h48;
mem[13198] = 8'hb9;
mem[13199] = 8'h5e;
mem[13200] = 8'h02;
mem[13201] = 8'h28;
mem[13202] = 8'h41;
mem[13203] = 8'h42;
mem[13204] = 8'h08;
mem[13205] = 8'hd9;
mem[13206] = 8'h62;
mem[13207] = 8'h02;
mem[13208] = 8'hd0;
mem[13209] = 8'hfe;
mem[13210] = 8'h68;
mem[13211] = 8'h09;
mem[13212] = 8'h08;
mem[13213] = 8'h49;
mem[13214] = 8'h38;
mem[13215] = 8'hd9;
mem[13216] = 8'h66;
mem[13217] = 8'h02;
mem[13218] = 8'hd0;
mem[13219] = 8'hfe;
mem[13220] = 8'hca;
mem[13221] = 8'hca;
mem[13222] = 8'h88;
mem[13223] = 8'h10;
mem[13224] = 8'he2;
mem[13225] = 8'ha2;
mem[13226] = 8'h06;
mem[13227] = 8'ha0;
mem[13228] = 8'h03;
mem[13229] = 8'ha9;
mem[13230] = 8'hff;
mem[13231] = 8'h48;
mem[13232] = 8'hb9;
mem[13233] = 8'h5e;
mem[13234] = 8'h02;
mem[13235] = 8'h28;
mem[13236] = 8'h41;
mem[13237] = 8'h42;
mem[13238] = 8'h08;
mem[13239] = 8'hd9;
mem[13240] = 8'h62;
mem[13241] = 8'h02;
mem[13242] = 8'hd0;
mem[13243] = 8'hfe;
mem[13244] = 8'h68;
mem[13245] = 8'h09;
mem[13246] = 8'h08;
mem[13247] = 8'h49;
mem[13248] = 8'h7d;
mem[13249] = 8'hd9;
mem[13250] = 8'h66;
mem[13251] = 8'h02;
mem[13252] = 8'hd0;
mem[13253] = 8'hfe;
mem[13254] = 8'hca;
mem[13255] = 8'hca;
mem[13256] = 8'h88;
mem[13257] = 8'h10;
mem[13258] = 8'he2;
mem[13259] = 8'ha0;
mem[13260] = 8'h03;
mem[13261] = 8'ha9;
mem[13262] = 8'h00;
mem[13263] = 8'h48;
mem[13264] = 8'hb9;
mem[13265] = 8'h5e;
mem[13266] = 8'h02;
mem[13267] = 8'h28;
mem[13268] = 8'h51;
mem[13269] = 8'h42;
mem[13270] = 8'h08;
mem[13271] = 8'hd9;
mem[13272] = 8'h62;
mem[13273] = 8'h02;
mem[13274] = 8'hd0;
mem[13275] = 8'hfe;
mem[13276] = 8'h68;
mem[13277] = 8'h09;
mem[13278] = 8'h08;
mem[13279] = 8'h49;
mem[13280] = 8'h38;
mem[13281] = 8'hd9;
mem[13282] = 8'h66;
mem[13283] = 8'h02;
mem[13284] = 8'hd0;
mem[13285] = 8'hfe;
mem[13286] = 8'h88;
mem[13287] = 8'h10;
mem[13288] = 8'he4;
mem[13289] = 8'ha0;
mem[13290] = 8'h03;
mem[13291] = 8'ha9;
mem[13292] = 8'hff;
mem[13293] = 8'h48;
mem[13294] = 8'hb9;
mem[13295] = 8'h5e;
mem[13296] = 8'h02;
mem[13297] = 8'h28;
mem[13298] = 8'h51;
mem[13299] = 8'h42;
mem[13300] = 8'h08;
mem[13301] = 8'hd9;
mem[13302] = 8'h62;
mem[13303] = 8'h02;
mem[13304] = 8'hd0;
mem[13305] = 8'hfe;
mem[13306] = 8'h68;
mem[13307] = 8'h09;
mem[13308] = 8'h08;
mem[13309] = 8'h49;
mem[13310] = 8'h7d;
mem[13311] = 8'hd9;
mem[13312] = 8'h66;
mem[13313] = 8'h02;
mem[13314] = 8'hd0;
mem[13315] = 8'hfe;
mem[13316] = 8'h88;
mem[13317] = 8'h10;
mem[13318] = 8'he4;
mem[13319] = 8'had;
mem[13320] = 8'h00;
mem[13321] = 8'h02;
mem[13322] = 8'hc9;
mem[13323] = 8'h27;
mem[13324] = 8'hd0;
mem[13325] = 8'hfe;
mem[13326] = 8'ha9;
mem[13327] = 8'h28;
mem[13328] = 8'h8d;
mem[13329] = 8'h00;
mem[13330] = 8'h02;
mem[13331] = 8'ha2;
mem[13332] = 8'h03;
mem[13333] = 8'hb5;
mem[13334] = 8'h18;
mem[13335] = 8'h8d;
mem[13336] = 8'h0f;
mem[13337] = 8'h02;
mem[13338] = 8'ha9;
mem[13339] = 8'h00;
mem[13340] = 8'h48;
mem[13341] = 8'hbd;
mem[13342] = 8'h56;
mem[13343] = 8'h02;
mem[13344] = 8'h28;
mem[13345] = 8'h20;
mem[13346] = 8'h0e;
mem[13347] = 8'h02;
mem[13348] = 8'h08;
mem[13349] = 8'hdd;
mem[13350] = 8'h62;
mem[13351] = 8'h02;
mem[13352] = 8'hd0;
mem[13353] = 8'hfe;
mem[13354] = 8'h68;
mem[13355] = 8'h09;
mem[13356] = 8'h08;
mem[13357] = 8'h49;
mem[13358] = 8'h38;
mem[13359] = 8'hdd;
mem[13360] = 8'h66;
mem[13361] = 8'h02;
mem[13362] = 8'hd0;
mem[13363] = 8'hfe;
mem[13364] = 8'hca;
mem[13365] = 8'h10;
mem[13366] = 8'hde;
mem[13367] = 8'ha2;
mem[13368] = 8'h03;
mem[13369] = 8'hb5;
mem[13370] = 8'h18;
mem[13371] = 8'h8d;
mem[13372] = 8'h0f;
mem[13373] = 8'h02;
mem[13374] = 8'ha9;
mem[13375] = 8'hff;
mem[13376] = 8'h48;
mem[13377] = 8'hbd;
mem[13378] = 8'h56;
mem[13379] = 8'h02;
mem[13380] = 8'h28;
mem[13381] = 8'h20;
mem[13382] = 8'h0e;
mem[13383] = 8'h02;
mem[13384] = 8'h08;
mem[13385] = 8'hdd;
mem[13386] = 8'h62;
mem[13387] = 8'h02;
mem[13388] = 8'hd0;
mem[13389] = 8'hfe;
mem[13390] = 8'h68;
mem[13391] = 8'h09;
mem[13392] = 8'h08;
mem[13393] = 8'h49;
mem[13394] = 8'h7d;
mem[13395] = 8'hdd;
mem[13396] = 8'h66;
mem[13397] = 8'h02;
mem[13398] = 8'hd0;
mem[13399] = 8'hfe;
mem[13400] = 8'hca;
mem[13401] = 8'h10;
mem[13402] = 8'hde;
mem[13403] = 8'ha2;
mem[13404] = 8'h03;
mem[13405] = 8'hb5;
mem[13406] = 8'h18;
mem[13407] = 8'h85;
mem[13408] = 8'h0c;
mem[13409] = 8'ha9;
mem[13410] = 8'h00;
mem[13411] = 8'h48;
mem[13412] = 8'hbd;
mem[13413] = 8'h56;
mem[13414] = 8'h02;
mem[13415] = 8'h28;
mem[13416] = 8'h05;
mem[13417] = 8'h0c;
mem[13418] = 8'h08;
mem[13419] = 8'hdd;
mem[13420] = 8'h62;
mem[13421] = 8'h02;
mem[13422] = 8'hd0;
mem[13423] = 8'hfe;
mem[13424] = 8'h68;
mem[13425] = 8'h09;
mem[13426] = 8'h08;
mem[13427] = 8'h49;
mem[13428] = 8'h38;
mem[13429] = 8'hdd;
mem[13430] = 8'h66;
mem[13431] = 8'h02;
mem[13432] = 8'hd0;
mem[13433] = 8'hfe;
mem[13434] = 8'hca;
mem[13435] = 8'h10;
mem[13436] = 8'he0;
mem[13437] = 8'ha2;
mem[13438] = 8'h03;
mem[13439] = 8'hb5;
mem[13440] = 8'h18;
mem[13441] = 8'h85;
mem[13442] = 8'h0c;
mem[13443] = 8'ha9;
mem[13444] = 8'hff;
mem[13445] = 8'h48;
mem[13446] = 8'hbd;
mem[13447] = 8'h56;
mem[13448] = 8'h02;
mem[13449] = 8'h28;
mem[13450] = 8'h05;
mem[13451] = 8'h0c;
mem[13452] = 8'h08;
mem[13453] = 8'hdd;
mem[13454] = 8'h62;
mem[13455] = 8'h02;
mem[13456] = 8'hd0;
mem[13457] = 8'hfe;
mem[13458] = 8'h68;
mem[13459] = 8'h09;
mem[13460] = 8'h08;
mem[13461] = 8'h49;
mem[13462] = 8'h7d;
mem[13463] = 8'hdd;
mem[13464] = 8'h66;
mem[13465] = 8'h02;
mem[13466] = 8'hd0;
mem[13467] = 8'hfe;
mem[13468] = 8'hca;
mem[13469] = 8'h10;
mem[13470] = 8'he0;
mem[13471] = 8'ha2;
mem[13472] = 8'h03;
mem[13473] = 8'hb5;
mem[13474] = 8'h18;
mem[13475] = 8'h8d;
mem[13476] = 8'h03;
mem[13477] = 8'h02;
mem[13478] = 8'ha9;
mem[13479] = 8'h00;
mem[13480] = 8'h48;
mem[13481] = 8'hbd;
mem[13482] = 8'h56;
mem[13483] = 8'h02;
mem[13484] = 8'h28;
mem[13485] = 8'h0d;
mem[13486] = 8'h03;
mem[13487] = 8'h02;
mem[13488] = 8'h08;
mem[13489] = 8'hdd;
mem[13490] = 8'h62;
mem[13491] = 8'h02;
mem[13492] = 8'hd0;
mem[13493] = 8'hfe;
mem[13494] = 8'h68;
mem[13495] = 8'h09;
mem[13496] = 8'h08;
mem[13497] = 8'h49;
mem[13498] = 8'h38;
mem[13499] = 8'hdd;
mem[13500] = 8'h66;
mem[13501] = 8'h02;
mem[13502] = 8'hd0;
mem[13503] = 8'hfe;
mem[13504] = 8'hca;
mem[13505] = 8'h10;
mem[13506] = 8'hde;
mem[13507] = 8'ha2;
mem[13508] = 8'h03;
mem[13509] = 8'hb5;
mem[13510] = 8'h18;
mem[13511] = 8'h8d;
mem[13512] = 8'h03;
mem[13513] = 8'h02;
mem[13514] = 8'ha9;
mem[13515] = 8'hff;
mem[13516] = 8'h48;
mem[13517] = 8'hbd;
mem[13518] = 8'h56;
mem[13519] = 8'h02;
mem[13520] = 8'h28;
mem[13521] = 8'h0d;
mem[13522] = 8'h03;
mem[13523] = 8'h02;
mem[13524] = 8'h08;
mem[13525] = 8'hdd;
mem[13526] = 8'h62;
mem[13527] = 8'h02;
mem[13528] = 8'hd0;
mem[13529] = 8'hfe;
mem[13530] = 8'h68;
mem[13531] = 8'h09;
mem[13532] = 8'h08;
mem[13533] = 8'h49;
mem[13534] = 8'h7d;
mem[13535] = 8'hdd;
mem[13536] = 8'h66;
mem[13537] = 8'h02;
mem[13538] = 8'hd0;
mem[13539] = 8'hfe;
mem[13540] = 8'hca;
mem[13541] = 8'h10;
mem[13542] = 8'h02;
mem[13543] = 8'ha2;
mem[13544] = 8'h03;
mem[13545] = 8'ha9;
mem[13546] = 8'h00;
mem[13547] = 8'h48;
mem[13548] = 8'hbd;
mem[13549] = 8'h56;
mem[13550] = 8'h02;
mem[13551] = 8'h28;
mem[13552] = 8'h15;
mem[13553] = 8'h18;
mem[13554] = 8'h08;
mem[13555] = 8'hdd;
mem[13556] = 8'h62;
mem[13557] = 8'h02;
mem[13558] = 8'hd0;
mem[13559] = 8'hfe;
mem[13560] = 8'h68;
mem[13561] = 8'h09;
mem[13562] = 8'h08;
mem[13563] = 8'h49;
mem[13564] = 8'h38;
mem[13565] = 8'hdd;
mem[13566] = 8'h66;
mem[13567] = 8'h02;
mem[13568] = 8'hd0;
mem[13569] = 8'hfe;
mem[13570] = 8'hca;
mem[13571] = 8'h10;
mem[13572] = 8'he4;
mem[13573] = 8'ha2;
mem[13574] = 8'h03;
mem[13575] = 8'ha9;
mem[13576] = 8'hff;
mem[13577] = 8'h48;
mem[13578] = 8'hbd;
mem[13579] = 8'h56;
mem[13580] = 8'h02;
mem[13581] = 8'h28;
mem[13582] = 8'h15;
mem[13583] = 8'h18;
mem[13584] = 8'h08;
mem[13585] = 8'hdd;
mem[13586] = 8'h62;
mem[13587] = 8'h02;
mem[13588] = 8'hd0;
mem[13589] = 8'hfe;
mem[13590] = 8'h68;
mem[13591] = 8'h09;
mem[13592] = 8'h08;
mem[13593] = 8'h49;
mem[13594] = 8'h7d;
mem[13595] = 8'hdd;
mem[13596] = 8'h66;
mem[13597] = 8'h02;
mem[13598] = 8'hd0;
mem[13599] = 8'hfe;
mem[13600] = 8'hca;
mem[13601] = 8'h10;
mem[13602] = 8'he4;
mem[13603] = 8'ha2;
mem[13604] = 8'h03;
mem[13605] = 8'ha9;
mem[13606] = 8'h00;
mem[13607] = 8'h48;
mem[13608] = 8'hbd;
mem[13609] = 8'h56;
mem[13610] = 8'h02;
mem[13611] = 8'h28;
mem[13612] = 8'h1d;
mem[13613] = 8'h4a;
mem[13614] = 8'h02;
mem[13615] = 8'h08;
mem[13616] = 8'hdd;
mem[13617] = 8'h62;
mem[13618] = 8'h02;
mem[13619] = 8'hd0;
mem[13620] = 8'hfe;
mem[13621] = 8'h68;
mem[13622] = 8'h09;
mem[13623] = 8'h08;
mem[13624] = 8'h49;
mem[13625] = 8'h38;
mem[13626] = 8'hdd;
mem[13627] = 8'h66;
mem[13628] = 8'h02;
mem[13629] = 8'hd0;
mem[13630] = 8'hfe;
mem[13631] = 8'hca;
mem[13632] = 8'h10;
mem[13633] = 8'he3;
mem[13634] = 8'ha2;
mem[13635] = 8'h03;
mem[13636] = 8'ha9;
mem[13637] = 8'hff;
mem[13638] = 8'h48;
mem[13639] = 8'hbd;
mem[13640] = 8'h56;
mem[13641] = 8'h02;
mem[13642] = 8'h28;
mem[13643] = 8'h1d;
mem[13644] = 8'h4a;
mem[13645] = 8'h02;
mem[13646] = 8'h08;
mem[13647] = 8'hdd;
mem[13648] = 8'h62;
mem[13649] = 8'h02;
mem[13650] = 8'hd0;
mem[13651] = 8'hfe;
mem[13652] = 8'h68;
mem[13653] = 8'h09;
mem[13654] = 8'h08;
mem[13655] = 8'h49;
mem[13656] = 8'h7d;
mem[13657] = 8'hdd;
mem[13658] = 8'h66;
mem[13659] = 8'h02;
mem[13660] = 8'hd0;
mem[13661] = 8'hfe;
mem[13662] = 8'hca;
mem[13663] = 8'h10;
mem[13664] = 8'he3;
mem[13665] = 8'ha0;
mem[13666] = 8'h03;
mem[13667] = 8'ha9;
mem[13668] = 8'h00;
mem[13669] = 8'h48;
mem[13670] = 8'hb9;
mem[13671] = 8'h56;
mem[13672] = 8'h02;
mem[13673] = 8'h28;
mem[13674] = 8'h19;
mem[13675] = 8'h4a;
mem[13676] = 8'h02;
mem[13677] = 8'h08;
mem[13678] = 8'hd9;
mem[13679] = 8'h62;
mem[13680] = 8'h02;
mem[13681] = 8'hd0;
mem[13682] = 8'hfe;
mem[13683] = 8'h68;
mem[13684] = 8'h09;
mem[13685] = 8'h08;
mem[13686] = 8'h49;
mem[13687] = 8'h38;
mem[13688] = 8'hd9;
mem[13689] = 8'h66;
mem[13690] = 8'h02;
mem[13691] = 8'hd0;
mem[13692] = 8'hfe;
mem[13693] = 8'h88;
mem[13694] = 8'h10;
mem[13695] = 8'he3;
mem[13696] = 8'ha0;
mem[13697] = 8'h03;
mem[13698] = 8'ha9;
mem[13699] = 8'hff;
mem[13700] = 8'h48;
mem[13701] = 8'hb9;
mem[13702] = 8'h56;
mem[13703] = 8'h02;
mem[13704] = 8'h28;
mem[13705] = 8'h19;
mem[13706] = 8'h4a;
mem[13707] = 8'h02;
mem[13708] = 8'h08;
mem[13709] = 8'hd9;
mem[13710] = 8'h62;
mem[13711] = 8'h02;
mem[13712] = 8'hd0;
mem[13713] = 8'hfe;
mem[13714] = 8'h68;
mem[13715] = 8'h09;
mem[13716] = 8'h08;
mem[13717] = 8'h49;
mem[13718] = 8'h7d;
mem[13719] = 8'hd9;
mem[13720] = 8'h66;
mem[13721] = 8'h02;
mem[13722] = 8'hd0;
mem[13723] = 8'hfe;
mem[13724] = 8'h88;
mem[13725] = 8'h10;
mem[13726] = 8'he3;
mem[13727] = 8'ha2;
mem[13728] = 8'h06;
mem[13729] = 8'ha0;
mem[13730] = 8'h03;
mem[13731] = 8'ha9;
mem[13732] = 8'h00;
mem[13733] = 8'h48;
mem[13734] = 8'hb9;
mem[13735] = 8'h56;
mem[13736] = 8'h02;
mem[13737] = 8'h28;
mem[13738] = 8'h01;
mem[13739] = 8'h4a;
mem[13740] = 8'h08;
mem[13741] = 8'hd9;
mem[13742] = 8'h62;
mem[13743] = 8'h02;
mem[13744] = 8'hd0;
mem[13745] = 8'hfe;
mem[13746] = 8'h68;
mem[13747] = 8'h09;
mem[13748] = 8'h08;
mem[13749] = 8'h49;
mem[13750] = 8'h38;
mem[13751] = 8'hd9;
mem[13752] = 8'h66;
mem[13753] = 8'h02;
mem[13754] = 8'hd0;
mem[13755] = 8'hfe;
mem[13756] = 8'hca;
mem[13757] = 8'hca;
mem[13758] = 8'h88;
mem[13759] = 8'h10;
mem[13760] = 8'he2;
mem[13761] = 8'ha2;
mem[13762] = 8'h06;
mem[13763] = 8'ha0;
mem[13764] = 8'h03;
mem[13765] = 8'ha9;
mem[13766] = 8'hff;
mem[13767] = 8'h48;
mem[13768] = 8'hb9;
mem[13769] = 8'h56;
mem[13770] = 8'h02;
mem[13771] = 8'h28;
mem[13772] = 8'h01;
mem[13773] = 8'h4a;
mem[13774] = 8'h08;
mem[13775] = 8'hd9;
mem[13776] = 8'h62;
mem[13777] = 8'h02;
mem[13778] = 8'hd0;
mem[13779] = 8'hfe;
mem[13780] = 8'h68;
mem[13781] = 8'h09;
mem[13782] = 8'h08;
mem[13783] = 8'h49;
mem[13784] = 8'h7d;
mem[13785] = 8'hd9;
mem[13786] = 8'h66;
mem[13787] = 8'h02;
mem[13788] = 8'hd0;
mem[13789] = 8'hfe;
mem[13790] = 8'hca;
mem[13791] = 8'hca;
mem[13792] = 8'h88;
mem[13793] = 8'h10;
mem[13794] = 8'he2;
mem[13795] = 8'ha0;
mem[13796] = 8'h03;
mem[13797] = 8'ha9;
mem[13798] = 8'h00;
mem[13799] = 8'h48;
mem[13800] = 8'hb9;
mem[13801] = 8'h56;
mem[13802] = 8'h02;
mem[13803] = 8'h28;
mem[13804] = 8'h11;
mem[13805] = 8'h4a;
mem[13806] = 8'h08;
mem[13807] = 8'hd9;
mem[13808] = 8'h62;
mem[13809] = 8'h02;
mem[13810] = 8'hd0;
mem[13811] = 8'hfe;
mem[13812] = 8'h68;
mem[13813] = 8'h09;
mem[13814] = 8'h08;
mem[13815] = 8'h49;
mem[13816] = 8'h38;
mem[13817] = 8'hd9;
mem[13818] = 8'h66;
mem[13819] = 8'h02;
mem[13820] = 8'hd0;
mem[13821] = 8'hfe;
mem[13822] = 8'h88;
mem[13823] = 8'h10;
mem[13824] = 8'he4;
mem[13825] = 8'ha0;
mem[13826] = 8'h03;
mem[13827] = 8'ha9;
mem[13828] = 8'hff;
mem[13829] = 8'h48;
mem[13830] = 8'hb9;
mem[13831] = 8'h56;
mem[13832] = 8'h02;
mem[13833] = 8'h28;
mem[13834] = 8'h11;
mem[13835] = 8'h4a;
mem[13836] = 8'h08;
mem[13837] = 8'hd9;
mem[13838] = 8'h62;
mem[13839] = 8'h02;
mem[13840] = 8'hd0;
mem[13841] = 8'hfe;
mem[13842] = 8'h68;
mem[13843] = 8'h09;
mem[13844] = 8'h08;
mem[13845] = 8'h49;
mem[13846] = 8'h7d;
mem[13847] = 8'hd9;
mem[13848] = 8'h66;
mem[13849] = 8'h02;
mem[13850] = 8'hd0;
mem[13851] = 8'hfe;
mem[13852] = 8'h88;
mem[13853] = 8'h10;
mem[13854] = 8'he4;
mem[13855] = 8'h58;
mem[13856] = 8'had;
mem[13857] = 8'h00;
mem[13858] = 8'h02;
mem[13859] = 8'hc9;
mem[13860] = 8'h28;
mem[13861] = 8'hd0;
mem[13862] = 8'hfe;
mem[13863] = 8'ha9;
mem[13864] = 8'h29;
mem[13865] = 8'h8d;
mem[13866] = 8'h00;
mem[13867] = 8'h02;
mem[13868] = 8'hd8;
mem[13869] = 8'ha2;
mem[13870] = 8'h0e;
mem[13871] = 8'ha0;
mem[13872] = 8'hff;
mem[13873] = 8'ha9;
mem[13874] = 8'h00;
mem[13875] = 8'h85;
mem[13876] = 8'h0c;
mem[13877] = 8'h85;
mem[13878] = 8'h0d;
mem[13879] = 8'h85;
mem[13880] = 8'h0e;
mem[13881] = 8'h8d;
mem[13882] = 8'h03;
mem[13883] = 8'h02;
mem[13884] = 8'h85;
mem[13885] = 8'h0f;
mem[13886] = 8'h85;
mem[13887] = 8'h10;
mem[13888] = 8'ha9;
mem[13889] = 8'hff;
mem[13890] = 8'h85;
mem[13891] = 8'h12;
mem[13892] = 8'h8d;
mem[13893] = 8'h04;
mem[13894] = 8'h02;
mem[13895] = 8'ha9;
mem[13896] = 8'h02;
mem[13897] = 8'h85;
mem[13898] = 8'h11;
mem[13899] = 8'h18;
mem[13900] = 8'h20;
mem[13901] = 8'h97;
mem[13902] = 8'h36;
mem[13903] = 8'he6;
mem[13904] = 8'h0c;
mem[13905] = 8'he6;
mem[13906] = 8'h0f;
mem[13907] = 8'h08;
mem[13908] = 8'h08;
mem[13909] = 8'h68;
mem[13910] = 8'h29;
mem[13911] = 8'h82;
mem[13912] = 8'h28;
mem[13913] = 8'hd0;
mem[13914] = 8'h02;
mem[13915] = 8'he6;
mem[13916] = 8'h10;
mem[13917] = 8'h05;
mem[13918] = 8'h10;
mem[13919] = 8'h85;
mem[13920] = 8'h11;
mem[13921] = 8'h38;
mem[13922] = 8'h20;
mem[13923] = 8'h97;
mem[13924] = 8'h36;
mem[13925] = 8'hc6;
mem[13926] = 8'h0c;
mem[13927] = 8'he6;
mem[13928] = 8'h0d;
mem[13929] = 8'hd0;
mem[13930] = 8'he0;
mem[13931] = 8'ha9;
mem[13932] = 8'h00;
mem[13933] = 8'h85;
mem[13934] = 8'h10;
mem[13935] = 8'hee;
mem[13936] = 8'h03;
mem[13937] = 8'h02;
mem[13938] = 8'he6;
mem[13939] = 8'h0e;
mem[13940] = 8'h08;
mem[13941] = 8'h68;
mem[13942] = 8'h29;
mem[13943] = 8'h82;
mem[13944] = 8'h85;
mem[13945] = 8'h11;
mem[13946] = 8'hc6;
mem[13947] = 8'h12;
mem[13948] = 8'hce;
mem[13949] = 8'h04;
mem[13950] = 8'h02;
mem[13951] = 8'ha5;
mem[13952] = 8'h0e;
mem[13953] = 8'h85;
mem[13954] = 8'h0f;
mem[13955] = 8'hd0;
mem[13956] = 8'hc6;
mem[13957] = 8'had;
mem[13958] = 8'h00;
mem[13959] = 8'h02;
mem[13960] = 8'hc9;
mem[13961] = 8'h29;
mem[13962] = 8'hd0;
mem[13963] = 8'hfe;
mem[13964] = 8'ha9;
mem[13965] = 8'hf0;
mem[13966] = 8'h8d;
mem[13967] = 8'h00;
mem[13968] = 8'h02;
mem[13969] = 8'h4c;
mem[13970] = 8'h91;
mem[13971] = 8'h36;
mem[13972] = 8'h4c;
mem[13973] = 8'h00;
mem[13974] = 8'h04;
mem[13975] = 8'ha5;
mem[13976] = 8'h11;
mem[13977] = 8'h29;
mem[13978] = 8'h83;
mem[13979] = 8'h48;
mem[13980] = 8'ha5;
mem[13981] = 8'h0d;
mem[13982] = 8'h45;
mem[13983] = 8'h0e;
mem[13984] = 8'h30;
mem[13985] = 8'h0a;
mem[13986] = 8'ha5;
mem[13987] = 8'h0d;
mem[13988] = 8'h45;
mem[13989] = 8'h0f;
mem[13990] = 8'h10;
mem[13991] = 8'h04;
mem[13992] = 8'h68;
mem[13993] = 8'h09;
mem[13994] = 8'h40;
mem[13995] = 8'h48;
mem[13996] = 8'h68;
mem[13997] = 8'h85;
mem[13998] = 8'h11;
mem[13999] = 8'h08;
mem[14000] = 8'ha5;
mem[14001] = 8'h0d;
mem[14002] = 8'h65;
mem[14003] = 8'h0e;
mem[14004] = 8'h08;
mem[14005] = 8'hc5;
mem[14006] = 8'h0f;
mem[14007] = 8'hd0;
mem[14008] = 8'hfe;
mem[14009] = 8'h68;
mem[14010] = 8'h29;
mem[14011] = 8'hc3;
mem[14012] = 8'hc5;
mem[14013] = 8'h11;
mem[14014] = 8'hd0;
mem[14015] = 8'hfe;
mem[14016] = 8'h28;
mem[14017] = 8'h08;
mem[14018] = 8'ha5;
mem[14019] = 8'h0d;
mem[14020] = 8'he5;
mem[14021] = 8'h12;
mem[14022] = 8'h08;
mem[14023] = 8'hc5;
mem[14024] = 8'h0f;
mem[14025] = 8'hd0;
mem[14026] = 8'hfe;
mem[14027] = 8'h68;
mem[14028] = 8'h29;
mem[14029] = 8'hc3;
mem[14030] = 8'hc5;
mem[14031] = 8'h11;
mem[14032] = 8'hd0;
mem[14033] = 8'hfe;
mem[14034] = 8'h28;
mem[14035] = 8'h08;
mem[14036] = 8'ha5;
mem[14037] = 8'h0d;
mem[14038] = 8'h6d;
mem[14039] = 8'h03;
mem[14040] = 8'h02;
mem[14041] = 8'h08;
mem[14042] = 8'hc5;
mem[14043] = 8'h0f;
mem[14044] = 8'hd0;
mem[14045] = 8'hfe;
mem[14046] = 8'h68;
mem[14047] = 8'h29;
mem[14048] = 8'hc3;
mem[14049] = 8'hc5;
mem[14050] = 8'h11;
mem[14051] = 8'hd0;
mem[14052] = 8'hfe;
mem[14053] = 8'h28;
mem[14054] = 8'h08;
mem[14055] = 8'ha5;
mem[14056] = 8'h0d;
mem[14057] = 8'hed;
mem[14058] = 8'h04;
mem[14059] = 8'h02;
mem[14060] = 8'h08;
mem[14061] = 8'hc5;
mem[14062] = 8'h0f;
mem[14063] = 8'hd0;
mem[14064] = 8'hfe;
mem[14065] = 8'h68;
mem[14066] = 8'h29;
mem[14067] = 8'hc3;
mem[14068] = 8'hc5;
mem[14069] = 8'h11;
mem[14070] = 8'hd0;
mem[14071] = 8'hfe;
mem[14072] = 8'h28;
mem[14073] = 8'h08;
mem[14074] = 8'ha5;
mem[14075] = 8'h0e;
mem[14076] = 8'h8d;
mem[14077] = 8'h12;
mem[14078] = 8'h02;
mem[14079] = 8'ha5;
mem[14080] = 8'h0d;
mem[14081] = 8'h20;
mem[14082] = 8'h11;
mem[14083] = 8'h02;
mem[14084] = 8'h08;
mem[14085] = 8'hc5;
mem[14086] = 8'h0f;
mem[14087] = 8'hd0;
mem[14088] = 8'hfe;
mem[14089] = 8'h68;
mem[14090] = 8'h29;
mem[14091] = 8'hc3;
mem[14092] = 8'hc5;
mem[14093] = 8'h11;
mem[14094] = 8'hd0;
mem[14095] = 8'hfe;
mem[14096] = 8'h28;
mem[14097] = 8'h08;
mem[14098] = 8'ha5;
mem[14099] = 8'h12;
mem[14100] = 8'h8d;
mem[14101] = 8'h15;
mem[14102] = 8'h02;
mem[14103] = 8'ha5;
mem[14104] = 8'h0d;
mem[14105] = 8'h20;
mem[14106] = 8'h14;
mem[14107] = 8'h02;
mem[14108] = 8'h08;
mem[14109] = 8'hc5;
mem[14110] = 8'h0f;
mem[14111] = 8'hd0;
mem[14112] = 8'hfe;
mem[14113] = 8'h68;
mem[14114] = 8'h29;
mem[14115] = 8'hc3;
mem[14116] = 8'hc5;
mem[14117] = 8'h11;
mem[14118] = 8'hd0;
mem[14119] = 8'hfe;
mem[14120] = 8'h28;
mem[14121] = 8'h08;
mem[14122] = 8'ha5;
mem[14123] = 8'h0d;
mem[14124] = 8'h75;
mem[14125] = 8'h00;
mem[14126] = 8'h08;
mem[14127] = 8'hc5;
mem[14128] = 8'h0f;
mem[14129] = 8'hd0;
mem[14130] = 8'hfe;
mem[14131] = 8'h68;
mem[14132] = 8'h29;
mem[14133] = 8'hc3;
mem[14134] = 8'hc5;
mem[14135] = 8'h11;
mem[14136] = 8'hd0;
mem[14137] = 8'hfe;
mem[14138] = 8'h28;
mem[14139] = 8'h08;
mem[14140] = 8'ha5;
mem[14141] = 8'h0d;
mem[14142] = 8'hf5;
mem[14143] = 8'h04;
mem[14144] = 8'h08;
mem[14145] = 8'hc5;
mem[14146] = 8'h0f;
mem[14147] = 8'hd0;
mem[14148] = 8'hfe;
mem[14149] = 8'h68;
mem[14150] = 8'h29;
mem[14151] = 8'hc3;
mem[14152] = 8'hc5;
mem[14153] = 8'h11;
mem[14154] = 8'hd0;
mem[14155] = 8'hfe;
mem[14156] = 8'h28;
mem[14157] = 8'h08;
mem[14158] = 8'ha5;
mem[14159] = 8'h0d;
mem[14160] = 8'h7d;
mem[14161] = 8'hf5;
mem[14162] = 8'h01;
mem[14163] = 8'h08;
mem[14164] = 8'hc5;
mem[14165] = 8'h0f;
mem[14166] = 8'hd0;
mem[14167] = 8'hfe;
mem[14168] = 8'h68;
mem[14169] = 8'h29;
mem[14170] = 8'hc3;
mem[14171] = 8'hc5;
mem[14172] = 8'h11;
mem[14173] = 8'hd0;
mem[14174] = 8'hfe;
mem[14175] = 8'h28;
mem[14176] = 8'h08;
mem[14177] = 8'ha5;
mem[14178] = 8'h0d;
mem[14179] = 8'hfd;
mem[14180] = 8'hf6;
mem[14181] = 8'h01;
mem[14182] = 8'h08;
mem[14183] = 8'hc5;
mem[14184] = 8'h0f;
mem[14185] = 8'hd0;
mem[14186] = 8'hfe;
mem[14187] = 8'h68;
mem[14188] = 8'h29;
mem[14189] = 8'hc3;
mem[14190] = 8'hc5;
mem[14191] = 8'h11;
mem[14192] = 8'hd0;
mem[14193] = 8'hfe;
mem[14194] = 8'h28;
mem[14195] = 8'h08;
mem[14196] = 8'ha5;
mem[14197] = 8'h0d;
mem[14198] = 8'h79;
mem[14199] = 8'h04;
mem[14200] = 8'h01;
mem[14201] = 8'h08;
mem[14202] = 8'hc5;
mem[14203] = 8'h0f;
mem[14204] = 8'hd0;
mem[14205] = 8'hfe;
mem[14206] = 8'h68;
mem[14207] = 8'h29;
mem[14208] = 8'hc3;
mem[14209] = 8'hc5;
mem[14210] = 8'h11;
mem[14211] = 8'hd0;
mem[14212] = 8'hfe;
mem[14213] = 8'h28;
mem[14214] = 8'h08;
mem[14215] = 8'ha5;
mem[14216] = 8'h0d;
mem[14217] = 8'hf9;
mem[14218] = 8'h05;
mem[14219] = 8'h01;
mem[14220] = 8'h08;
mem[14221] = 8'hc5;
mem[14222] = 8'h0f;
mem[14223] = 8'hd0;
mem[14224] = 8'hfe;
mem[14225] = 8'h68;
mem[14226] = 8'h29;
mem[14227] = 8'hc3;
mem[14228] = 8'hc5;
mem[14229] = 8'h11;
mem[14230] = 8'hd0;
mem[14231] = 8'hfe;
mem[14232] = 8'h28;
mem[14233] = 8'h08;
mem[14234] = 8'ha5;
mem[14235] = 8'h0d;
mem[14236] = 8'h61;
mem[14237] = 8'h44;
mem[14238] = 8'h08;
mem[14239] = 8'hc5;
mem[14240] = 8'h0f;
mem[14241] = 8'hd0;
mem[14242] = 8'hfe;
mem[14243] = 8'h68;
mem[14244] = 8'h29;
mem[14245] = 8'hc3;
mem[14246] = 8'hc5;
mem[14247] = 8'h11;
mem[14248] = 8'hd0;
mem[14249] = 8'hfe;
mem[14250] = 8'h28;
mem[14251] = 8'h08;
mem[14252] = 8'ha5;
mem[14253] = 8'h0d;
mem[14254] = 8'he1;
mem[14255] = 8'h46;
mem[14256] = 8'h08;
mem[14257] = 8'hc5;
mem[14258] = 8'h0f;
mem[14259] = 8'hd0;
mem[14260] = 8'hfe;
mem[14261] = 8'h68;
mem[14262] = 8'h29;
mem[14263] = 8'hc3;
mem[14264] = 8'hc5;
mem[14265] = 8'h11;
mem[14266] = 8'hd0;
mem[14267] = 8'hfe;
mem[14268] = 8'h28;
mem[14269] = 8'h08;
mem[14270] = 8'ha5;
mem[14271] = 8'h0d;
mem[14272] = 8'h71;
mem[14273] = 8'h56;
mem[14274] = 8'h08;
mem[14275] = 8'hc5;
mem[14276] = 8'h0f;
mem[14277] = 8'hd0;
mem[14278] = 8'hfe;
mem[14279] = 8'h68;
mem[14280] = 8'h29;
mem[14281] = 8'hc3;
mem[14282] = 8'hc5;
mem[14283] = 8'h11;
mem[14284] = 8'hd0;
mem[14285] = 8'hfe;
mem[14286] = 8'h28;
mem[14287] = 8'h08;
mem[14288] = 8'ha5;
mem[14289] = 8'h0d;
mem[14290] = 8'hf1;
mem[14291] = 8'h58;
mem[14292] = 8'h08;
mem[14293] = 8'hc5;
mem[14294] = 8'h0f;
mem[14295] = 8'hd0;
mem[14296] = 8'hfe;
mem[14297] = 8'h68;
mem[14298] = 8'h29;
mem[14299] = 8'hc3;
mem[14300] = 8'hc5;
mem[14301] = 8'h11;
mem[14302] = 8'hd0;
mem[14303] = 8'hfe;
mem[14304] = 8'h28;
mem[14305] = 8'h60;
mem[14306] = 8'h88;
mem[14307] = 8'h88;
mem[14308] = 8'h08;
mem[14309] = 8'h88;
mem[14310] = 8'h88;
mem[14311] = 8'h88;
mem[14312] = 8'h28;
mem[14313] = 8'hb0;
mem[14314] = 8'hfe;
mem[14315] = 8'h70;
mem[14316] = 8'hfe;
mem[14317] = 8'h30;
mem[14318] = 8'hfe;
mem[14319] = 8'hf0;
mem[14320] = 8'hfe;
mem[14321] = 8'hc9;
mem[14322] = 8'h46;
mem[14323] = 8'hd0;
mem[14324] = 8'hfe;
mem[14325] = 8'he0;
mem[14326] = 8'h41;
mem[14327] = 8'hd0;
mem[14328] = 8'hfe;
mem[14329] = 8'hc0;
mem[14330] = 8'h4f;
mem[14331] = 8'hd0;
mem[14332] = 8'hfe;
mem[14333] = 8'h48;
mem[14334] = 8'h8a;
mem[14335] = 8'h48;
mem[14336] = 8'hba;
mem[14337] = 8'he0;
mem[14338] = 8'hfd;
mem[14339] = 8'hd0;
mem[14340] = 8'hfe;
mem[14341] = 8'h68;
mem[14342] = 8'haa;
mem[14343] = 8'ha9;
mem[14344] = 8'hff;
mem[14345] = 8'h48;
mem[14346] = 8'h28;
mem[14347] = 8'h68;
mem[14348] = 8'he8;
mem[14349] = 8'h49;
mem[14350] = 8'haa;
mem[14351] = 8'h4c;
mem[14352] = 8'h53;
mem[14353] = 8'h09;
mem[14354] = 8'h1b;
mem[14355] = 8'h38;
mem[14356] = 8'ha8;
mem[14357] = 8'h09;
mem[14358] = 8'h4c;
mem[14359] = 8'h16;
mem[14360] = 8'h38;
mem[14361] = 8'h88;
mem[14362] = 8'h88;
mem[14363] = 8'h08;
mem[14364] = 8'h88;
mem[14365] = 8'h88;
mem[14366] = 8'h88;
mem[14367] = 8'h28;
mem[14368] = 8'hb0;
mem[14369] = 8'hfe;
mem[14370] = 8'h70;
mem[14371] = 8'hfe;
mem[14372] = 8'h30;
mem[14373] = 8'hfe;
mem[14374] = 8'hf0;
mem[14375] = 8'hfe;
mem[14376] = 8'hc9;
mem[14377] = 8'h49;
mem[14378] = 8'hd0;
mem[14379] = 8'hfe;
mem[14380] = 8'he0;
mem[14381] = 8'h4e;
mem[14382] = 8'hd0;
mem[14383] = 8'hfe;
mem[14384] = 8'hc0;
mem[14385] = 8'h41;
mem[14386] = 8'hd0;
mem[14387] = 8'hfe;
mem[14388] = 8'h48;
mem[14389] = 8'h8a;
mem[14390] = 8'h48;
mem[14391] = 8'hba;
mem[14392] = 8'he0;
mem[14393] = 8'hfd;
mem[14394] = 8'hd0;
mem[14395] = 8'hfe;
mem[14396] = 8'h68;
mem[14397] = 8'haa;
mem[14398] = 8'ha9;
mem[14399] = 8'hff;
mem[14400] = 8'h48;
mem[14401] = 8'h28;
mem[14402] = 8'h68;
mem[14403] = 8'he8;
mem[14404] = 8'h49;
mem[14405] = 8'haa;
mem[14406] = 8'h6c;
mem[14407] = 8'h14;
mem[14408] = 8'h38;
mem[14409] = 8'h4c;
mem[14410] = 8'h49;
mem[14411] = 8'h38;
mem[14412] = 8'h88;
mem[14413] = 8'h88;
mem[14414] = 8'h08;
mem[14415] = 8'h88;
mem[14416] = 8'h88;
mem[14417] = 8'h88;
mem[14418] = 8'h28;
mem[14419] = 8'hb0;
mem[14420] = 8'hfe;
mem[14421] = 8'h70;
mem[14422] = 8'hfe;
mem[14423] = 8'h30;
mem[14424] = 8'hfe;
mem[14425] = 8'hf0;
mem[14426] = 8'hfe;
mem[14427] = 8'hc9;
mem[14428] = 8'h4a;
mem[14429] = 8'hd0;
mem[14430] = 8'hfe;
mem[14431] = 8'he0;
mem[14432] = 8'h53;
mem[14433] = 8'hd0;
mem[14434] = 8'hfe;
mem[14435] = 8'hc0;
mem[14436] = 8'h4f;
mem[14437] = 8'hd0;
mem[14438] = 8'hfe;
mem[14439] = 8'h48;
mem[14440] = 8'h8a;
mem[14441] = 8'h48;
mem[14442] = 8'hba;
mem[14443] = 8'he0;
mem[14444] = 8'hfb;
mem[14445] = 8'hd0;
mem[14446] = 8'hfe;
mem[14447] = 8'had;
mem[14448] = 8'hff;
mem[14449] = 8'h01;
mem[14450] = 8'hc9;
mem[14451] = 8'h09;
mem[14452] = 8'hd0;
mem[14453] = 8'hfe;
mem[14454] = 8'had;
mem[14455] = 8'hfe;
mem[14456] = 8'h01;
mem[14457] = 8'hc9;
mem[14458] = 8'hde;
mem[14459] = 8'hd0;
mem[14460] = 8'hfe;
mem[14461] = 8'ha9;
mem[14462] = 8'hff;
mem[14463] = 8'h48;
mem[14464] = 8'h28;
mem[14465] = 8'h68;
mem[14466] = 8'haa;
mem[14467] = 8'h68;
mem[14468] = 8'he8;
mem[14469] = 8'h49;
mem[14470] = 8'haa;
mem[14471] = 8'h60;
mem[14472] = 8'h4c;
mem[14473] = 8'h88;
mem[14474] = 8'h38;
mem[14475] = 8'h4c;
mem[14476] = 8'h8b;
mem[14477] = 8'h38;
mem[14478] = 8'h4c;
mem[14479] = 8'h8e;
mem[14480] = 8'h38;
mem[14481] = 8'h88;
mem[14482] = 8'h88;
mem[14483] = 8'h08;
mem[14484] = 8'h88;
mem[14485] = 8'h88;
mem[14486] = 8'h88;
mem[14487] = 8'hc9;
mem[14488] = 8'h42;
mem[14489] = 8'hd0;
mem[14490] = 8'hfe;
mem[14491] = 8'he0;
mem[14492] = 8'h52;
mem[14493] = 8'hd0;
mem[14494] = 8'hfe;
mem[14495] = 8'hc0;
mem[14496] = 8'h48;
mem[14497] = 8'hd0;
mem[14498] = 8'hfe;
mem[14499] = 8'h85;
mem[14500] = 8'h0a;
mem[14501] = 8'h86;
mem[14502] = 8'h0b;
mem[14503] = 8'hba;
mem[14504] = 8'hbd;
mem[14505] = 8'h02;
mem[14506] = 8'h01;
mem[14507] = 8'h09;
mem[14508] = 8'h08;
mem[14509] = 8'hc9;
mem[14510] = 8'h38;
mem[14511] = 8'hd0;
mem[14512] = 8'hfe;
mem[14513] = 8'h68;
mem[14514] = 8'hc9;
mem[14515] = 8'h34;
mem[14516] = 8'hd0;
mem[14517] = 8'hfe;
mem[14518] = 8'hba;
mem[14519] = 8'he0;
mem[14520] = 8'hfc;
mem[14521] = 8'hd0;
mem[14522] = 8'hfe;
mem[14523] = 8'had;
mem[14524] = 8'hff;
mem[14525] = 8'h01;
mem[14526] = 8'hc9;
mem[14527] = 8'h0a;
mem[14528] = 8'hd0;
mem[14529] = 8'hfe;
mem[14530] = 8'had;
mem[14531] = 8'hfe;
mem[14532] = 8'h01;
mem[14533] = 8'hc9;
mem[14534] = 8'h15;
mem[14535] = 8'hd0;
mem[14536] = 8'hfe;
mem[14537] = 8'ha9;
mem[14538] = 8'hff;
mem[14539] = 8'h48;
mem[14540] = 8'h28;
mem[14541] = 8'ha6;
mem[14542] = 8'h0b;
mem[14543] = 8'he8;
mem[14544] = 8'ha5;
mem[14545] = 8'h0a;
mem[14546] = 8'h49;
mem[14547] = 8'haa;
mem[14548] = 8'h40;
mem[14549] = 8'h4c;
mem[14550] = 8'hd5;
mem[14551] = 8'h38;
mem[14552] = 8'hc3;
mem[14553] = 8'h82;
mem[14554] = 8'h41;
mem[14555] = 8'h00;
mem[14556] = 8'h7f;
mem[14557] = 8'h00;
mem[14558] = 8'h1f;
mem[14559] = 8'h71;
mem[14560] = 8'h80;
mem[14561] = 8'h0f;
mem[14562] = 8'hff;
mem[14563] = 8'h7f;
mem[14564] = 8'h80;
mem[14565] = 8'hff;
mem[14566] = 8'h0f;
mem[14567] = 8'h8f;
mem[14568] = 8'h8f;
mem[14569] = 8'h17;
mem[14570] = 8'h02;
mem[14571] = 8'h18;
mem[14572] = 8'h02;
mem[14573] = 8'h19;
mem[14574] = 8'h02;
mem[14575] = 8'h1a;
mem[14576] = 8'h02;
mem[14577] = 8'h1b;
mem[14578] = 8'h02;
mem[14579] = 8'h1f;
mem[14580] = 8'h01;
mem[14581] = 8'h03;
mem[14582] = 8'h02;
mem[14583] = 8'h04;
mem[14584] = 8'h02;
mem[14585] = 8'h05;
mem[14586] = 8'h02;
mem[14587] = 8'h06;
mem[14588] = 8'h02;
mem[14589] = 8'h0b;
mem[14590] = 8'h01;
mem[14591] = 8'h4e;
mem[14592] = 8'h02;
mem[14593] = 8'h4f;
mem[14594] = 8'h02;
mem[14595] = 8'h50;
mem[14596] = 8'h02;
mem[14597] = 8'h51;
mem[14598] = 8'h02;
mem[14599] = 8'h52;
mem[14600] = 8'h02;
mem[14601] = 8'h53;
mem[14602] = 8'h02;
mem[14603] = 8'h54;
mem[14604] = 8'h02;
mem[14605] = 8'h55;
mem[14606] = 8'h02;
mem[14607] = 8'h4a;
mem[14608] = 8'h02;
mem[14609] = 8'h4b;
mem[14610] = 8'h02;
mem[14611] = 8'h4c;
mem[14612] = 8'h02;
mem[14613] = 8'h4d;
mem[14614] = 8'h02;
mem[14615] = 8'h03;
mem[14616] = 8'h02;
mem[14617] = 8'h04;
mem[14618] = 8'h02;
mem[14619] = 8'h04;
mem[14620] = 8'h01;
mem[14621] = 8'h05;
mem[14622] = 8'h01;
mem[14623] = 8'h29;
mem[14624] = 8'h00;
mem[14625] = 8'h60;
mem[14626] = 8'h49;
mem[14627] = 8'h00;
mem[14628] = 8'h60;
mem[14629] = 8'h09;
mem[14630] = 8'h00;
mem[14631] = 8'h60;
mem[14632] = 8'h69;
mem[14633] = 8'h00;
mem[14634] = 8'h60;
mem[14635] = 8'he9;
mem[14636] = 8'h00;
mem[14637] = 8'h60;
mem[14638] = 8'hc3;
mem[14639] = 8'h82;
mem[14640] = 8'h41;
mem[14641] = 8'h00;
mem[14642] = 8'h7f;
mem[14643] = 8'h80;
mem[14644] = 8'h80;
mem[14645] = 8'h00;
mem[14646] = 8'h02;
mem[14647] = 8'h86;
mem[14648] = 8'h04;
mem[14649] = 8'h82;
mem[14650] = 8'h00;
mem[14651] = 8'h87;
mem[14652] = 8'h05;
mem[14653] = 8'h83;
mem[14654] = 8'h01;
mem[14655] = 8'h61;
mem[14656] = 8'h41;
mem[14657] = 8'h20;
mem[14658] = 8'h00;
mem[14659] = 8'he1;
mem[14660] = 8'hc1;
mem[14661] = 8'ha0;
mem[14662] = 8'h80;
mem[14663] = 8'h81;
mem[14664] = 8'h01;
mem[14665] = 8'h80;
mem[14666] = 8'h02;
mem[14667] = 8'h81;
mem[14668] = 8'h01;
mem[14669] = 8'h80;
mem[14670] = 8'h00;
mem[14671] = 8'h01;
mem[14672] = 8'h00;
mem[14673] = 8'h01;
mem[14674] = 8'h02;
mem[14675] = 8'h81;
mem[14676] = 8'h80;
mem[14677] = 8'h81;
mem[14678] = 8'h80;
mem[14679] = 8'h7f;
mem[14680] = 8'h80;
mem[14681] = 8'hff;
mem[14682] = 8'h00;
mem[14683] = 8'h01;
mem[14684] = 8'h00;
mem[14685] = 8'h80;
mem[14686] = 8'h80;
mem[14687] = 8'h02;
mem[14688] = 8'h00;
mem[14689] = 8'h00;
mem[14690] = 8'h1f;
mem[14691] = 8'h71;
mem[14692] = 8'h80;
mem[14693] = 8'h0f;
mem[14694] = 8'hff;
mem[14695] = 8'h7f;
mem[14696] = 8'h80;
mem[14697] = 8'hff;
mem[14698] = 8'h0f;
mem[14699] = 8'h8f;
mem[14700] = 8'h8f;
mem[14701] = 8'h00;
mem[14702] = 8'hf1;
mem[14703] = 8'h1f;
mem[14704] = 8'h00;
mem[14705] = 8'hf0;
mem[14706] = 8'hff;
mem[14707] = 8'hff;
mem[14708] = 8'hff;
mem[14709] = 8'hff;
mem[14710] = 8'hf0;
mem[14711] = 8'hf0;
mem[14712] = 8'h0f;
mem[14713] = 8'h00;
mem[14714] = 8'hff;
mem[14715] = 8'h7f;
mem[14716] = 8'h80;
mem[14717] = 8'h02;
mem[14718] = 8'h80;
mem[14719] = 8'h00;
mem[14720] = 8'h80;
mem[14721] = 8'h8b;
mem[14722] = 8'h38;
mem[14723] = 8'h8e;
mem[14724] = 8'h38;
mem[14725] = 8'h93;
mem[14726] = 8'h38;
mem[14727] = 8'h00;
mem[14728] = 8'h00;
mem[14729] = 8'h00;
mem[14730] = 8'h00;
mem[14731] = 8'h00;
mem[14732] = 8'h00;
mem[14733] = 8'h00;
mem[14734] = 8'h00;
mem[14735] = 8'h00;
mem[14736] = 8'h00;
mem[14737] = 8'h00;
mem[14738] = 8'h00;
mem[14739] = 8'h00;
mem[14740] = 8'h00;
mem[14741] = 8'h00;
mem[14742] = 8'h00;
mem[14743] = 8'h00;
mem[14744] = 8'h00;
mem[14745] = 8'h00;
mem[14746] = 8'h00;
mem[14747] = 8'h00;
mem[14748] = 8'h00;
mem[14749] = 8'h00;
mem[14750] = 8'h00;
mem[14751] = 8'h00;
mem[14752] = 8'h00;
mem[14753] = 8'h00;
mem[14754] = 8'h00;
mem[14755] = 8'h00;
mem[14756] = 8'h00;
mem[14757] = 8'h00;
mem[14758] = 8'h00;
mem[14759] = 8'h00;
mem[14760] = 8'h00;
mem[14761] = 8'h00;
mem[14762] = 8'h00;
mem[14763] = 8'h00;
mem[14764] = 8'h00;
mem[14765] = 8'h00;
mem[14766] = 8'h00;
mem[14767] = 8'h00;
mem[14768] = 8'h00;
mem[14769] = 8'h00;
mem[14770] = 8'h00;
mem[14771] = 8'h00;
mem[14772] = 8'h00;
mem[14773] = 8'h00;
mem[14774] = 8'h00;
mem[14775] = 8'h00;
mem[14776] = 8'h00;
mem[14777] = 8'h00;
mem[14778] = 8'h00;
mem[14779] = 8'h00;
mem[14780] = 8'h00;
mem[14781] = 8'h00;
mem[14782] = 8'h00;
mem[14783] = 8'h00;
mem[14784] = 8'h00;
mem[14785] = 8'h00;
mem[14786] = 8'h00;
mem[14787] = 8'h00;
mem[14788] = 8'h00;
mem[14789] = 8'h00;
mem[14790] = 8'h00;
mem[14791] = 8'h00;
mem[14792] = 8'h00;
mem[14793] = 8'h00;
mem[14794] = 8'h00;
mem[14795] = 8'h00;
mem[14796] = 8'h00;
mem[14797] = 8'h00;
mem[14798] = 8'h00;
mem[14799] = 8'h00;
mem[14800] = 8'h00;
mem[14801] = 8'h00;
mem[14802] = 8'h00;
mem[14803] = 8'h00;
mem[14804] = 8'h00;
mem[14805] = 8'h00;
mem[14806] = 8'h00;
mem[14807] = 8'h00;
mem[14808] = 8'h00;
mem[14809] = 8'h00;
mem[14810] = 8'h00;
mem[14811] = 8'h00;
mem[14812] = 8'h00;
mem[14813] = 8'h00;
mem[14814] = 8'h00;
mem[14815] = 8'h00;
mem[14816] = 8'h00;
mem[14817] = 8'h00;
mem[14818] = 8'h00;
mem[14819] = 8'h00;
mem[14820] = 8'h00;
mem[14821] = 8'h00;
mem[14822] = 8'h00;
mem[14823] = 8'h00;
mem[14824] = 8'h00;
mem[14825] = 8'h00;
mem[14826] = 8'h00;
mem[14827] = 8'h00;
mem[14828] = 8'h00;
mem[14829] = 8'h00;
mem[14830] = 8'h00;
mem[14831] = 8'h00;
mem[14832] = 8'h00;
mem[14833] = 8'h00;
mem[14834] = 8'h00;
mem[14835] = 8'h00;
mem[14836] = 8'h00;
mem[14837] = 8'h00;
mem[14838] = 8'h00;
mem[14839] = 8'h00;
mem[14840] = 8'h00;
mem[14841] = 8'h00;
mem[14842] = 8'h00;
mem[14843] = 8'h00;
mem[14844] = 8'h00;
mem[14845] = 8'h00;
mem[14846] = 8'h00;
mem[14847] = 8'h00;
mem[14848] = 8'h00;
mem[14849] = 8'h00;
mem[14850] = 8'h00;
mem[14851] = 8'h00;
mem[14852] = 8'h00;
mem[14853] = 8'h00;
mem[14854] = 8'h00;
mem[14855] = 8'h00;
mem[14856] = 8'h00;
mem[14857] = 8'h00;
mem[14858] = 8'h00;
mem[14859] = 8'h00;
mem[14860] = 8'h00;
mem[14861] = 8'h00;
mem[14862] = 8'h00;
mem[14863] = 8'h00;
mem[14864] = 8'h00;
mem[14865] = 8'h00;
mem[14866] = 8'h00;
mem[14867] = 8'h00;
mem[14868] = 8'h00;
mem[14869] = 8'h00;
mem[14870] = 8'h00;
mem[14871] = 8'h00;
mem[14872] = 8'h00;
mem[14873] = 8'h00;
mem[14874] = 8'h00;
mem[14875] = 8'h00;
mem[14876] = 8'h00;
mem[14877] = 8'h00;
mem[14878] = 8'h00;
mem[14879] = 8'h00;
mem[14880] = 8'h00;
mem[14881] = 8'h00;
mem[14882] = 8'h00;
mem[14883] = 8'h00;
mem[14884] = 8'h00;
mem[14885] = 8'h00;
mem[14886] = 8'h00;
mem[14887] = 8'h00;
mem[14888] = 8'h00;
mem[14889] = 8'h00;
mem[14890] = 8'h00;
mem[14891] = 8'h00;
mem[14892] = 8'h00;
mem[14893] = 8'h00;
mem[14894] = 8'h00;
mem[14895] = 8'h00;
mem[14896] = 8'h00;
mem[14897] = 8'h00;
mem[14898] = 8'h00;
mem[14899] = 8'h00;
mem[14900] = 8'h00;
mem[14901] = 8'h00;
mem[14902] = 8'h00;
mem[14903] = 8'h00;
mem[14904] = 8'h00;
mem[14905] = 8'h00;
mem[14906] = 8'h00;
mem[14907] = 8'h00;
mem[14908] = 8'h00;
mem[14909] = 8'h00;
mem[14910] = 8'h00;
mem[14911] = 8'h00;
mem[14912] = 8'h00;
mem[14913] = 8'h00;
mem[14914] = 8'h00;
mem[14915] = 8'h00;
mem[14916] = 8'h00;
mem[14917] = 8'h00;
mem[14918] = 8'h00;
mem[14919] = 8'h00;
mem[14920] = 8'h00;
mem[14921] = 8'h00;
mem[14922] = 8'h00;
mem[14923] = 8'h00;
mem[14924] = 8'h00;
mem[14925] = 8'h00;
mem[14926] = 8'h00;
mem[14927] = 8'h00;
mem[14928] = 8'h00;
mem[14929] = 8'h00;
mem[14930] = 8'h00;
mem[14931] = 8'h00;
mem[14932] = 8'h00;
mem[14933] = 8'h00;
mem[14934] = 8'h00;
mem[14935] = 8'h00;
mem[14936] = 8'h00;
mem[14937] = 8'h00;
mem[14938] = 8'h00;
mem[14939] = 8'h00;
mem[14940] = 8'h00;
mem[14941] = 8'h00;
mem[14942] = 8'h00;
mem[14943] = 8'h00;
mem[14944] = 8'h00;
mem[14945] = 8'h00;
mem[14946] = 8'h00;
mem[14947] = 8'h00;
mem[14948] = 8'h00;
mem[14949] = 8'h00;
mem[14950] = 8'h00;
mem[14951] = 8'h00;
mem[14952] = 8'h00;
mem[14953] = 8'h00;
mem[14954] = 8'h00;
mem[14955] = 8'h00;
mem[14956] = 8'h00;
mem[14957] = 8'h00;
mem[14958] = 8'h00;
mem[14959] = 8'h00;
mem[14960] = 8'h00;
mem[14961] = 8'h00;
mem[14962] = 8'h00;
mem[14963] = 8'h00;
mem[14964] = 8'h00;
mem[14965] = 8'h00;
mem[14966] = 8'h00;
mem[14967] = 8'h00;
mem[14968] = 8'h00;
mem[14969] = 8'h00;
mem[14970] = 8'h00;
mem[14971] = 8'h00;
mem[14972] = 8'h00;
mem[14973] = 8'h00;
mem[14974] = 8'h00;
mem[14975] = 8'h00;
mem[14976] = 8'h00;
mem[14977] = 8'h00;
mem[14978] = 8'h00;
mem[14979] = 8'h00;
mem[14980] = 8'h00;
mem[14981] = 8'h00;
mem[14982] = 8'h00;
mem[14983] = 8'h00;
mem[14984] = 8'h00;
mem[14985] = 8'h00;
mem[14986] = 8'h00;
mem[14987] = 8'h00;
mem[14988] = 8'h00;
mem[14989] = 8'h00;
mem[14990] = 8'h00;
mem[14991] = 8'h00;
mem[14992] = 8'h00;
mem[14993] = 8'h00;
mem[14994] = 8'h00;
mem[14995] = 8'h00;
mem[14996] = 8'h00;
mem[14997] = 8'h00;
mem[14998] = 8'h00;
mem[14999] = 8'h00;
mem[15000] = 8'h00;
mem[15001] = 8'h00;
mem[15002] = 8'h00;
mem[15003] = 8'h00;
mem[15004] = 8'h00;
mem[15005] = 8'h00;
mem[15006] = 8'h00;
mem[15007] = 8'h00;
mem[15008] = 8'h00;
mem[15009] = 8'h00;
mem[15010] = 8'h00;
mem[15011] = 8'h00;
mem[15012] = 8'h00;
mem[15013] = 8'h00;
mem[15014] = 8'h00;
mem[15015] = 8'h00;
mem[15016] = 8'h00;
mem[15017] = 8'h00;
mem[15018] = 8'h00;
mem[15019] = 8'h00;
mem[15020] = 8'h00;
mem[15021] = 8'h00;
mem[15022] = 8'h00;
mem[15023] = 8'h00;
mem[15024] = 8'h00;
mem[15025] = 8'h00;
mem[15026] = 8'h00;
mem[15027] = 8'h00;
mem[15028] = 8'h00;
mem[15029] = 8'h00;
mem[15030] = 8'h00;
mem[15031] = 8'h00;
mem[15032] = 8'h00;
mem[15033] = 8'h00;
mem[15034] = 8'h00;
mem[15035] = 8'h00;
mem[15036] = 8'h00;
mem[15037] = 8'h00;
mem[15038] = 8'h00;
mem[15039] = 8'h00;
mem[15040] = 8'h00;
mem[15041] = 8'h00;
mem[15042] = 8'h00;
mem[15043] = 8'h00;
mem[15044] = 8'h00;
mem[15045] = 8'h00;
mem[15046] = 8'h00;
mem[15047] = 8'h00;
mem[15048] = 8'h00;
mem[15049] = 8'h00;
mem[15050] = 8'h00;
mem[15051] = 8'h00;
mem[15052] = 8'h00;
mem[15053] = 8'h00;
mem[15054] = 8'h00;
mem[15055] = 8'h00;
mem[15056] = 8'h00;
mem[15057] = 8'h00;
mem[15058] = 8'h00;
mem[15059] = 8'h00;
mem[15060] = 8'h00;
mem[15061] = 8'h00;
mem[15062] = 8'h00;
mem[15063] = 8'h00;
mem[15064] = 8'h00;
mem[15065] = 8'h00;
mem[15066] = 8'h00;
mem[15067] = 8'h00;
mem[15068] = 8'h00;
mem[15069] = 8'h00;
mem[15070] = 8'h00;
mem[15071] = 8'h00;
mem[15072] = 8'h00;
mem[15073] = 8'h00;
mem[15074] = 8'h00;
mem[15075] = 8'h00;
mem[15076] = 8'h00;
mem[15077] = 8'h00;
mem[15078] = 8'h00;
mem[15079] = 8'h00;
mem[15080] = 8'h00;
mem[15081] = 8'h00;
mem[15082] = 8'h00;
mem[15083] = 8'h00;
mem[15084] = 8'h00;
mem[15085] = 8'h00;
mem[15086] = 8'h00;
mem[15087] = 8'h00;
mem[15088] = 8'h00;
mem[15089] = 8'h00;
mem[15090] = 8'h00;
mem[15091] = 8'h00;
mem[15092] = 8'h00;
mem[15093] = 8'h00;
mem[15094] = 8'h00;
mem[15095] = 8'h00;
mem[15096] = 8'h00;
mem[15097] = 8'h00;
mem[15098] = 8'h00;
mem[15099] = 8'h00;
mem[15100] = 8'h00;
mem[15101] = 8'h00;
mem[15102] = 8'h00;
mem[15103] = 8'h00;
mem[15104] = 8'h00;
mem[15105] = 8'h00;
mem[15106] = 8'h00;
mem[15107] = 8'h00;
mem[15108] = 8'h00;
mem[15109] = 8'h00;
mem[15110] = 8'h00;
mem[15111] = 8'h00;
mem[15112] = 8'h00;
mem[15113] = 8'h00;
mem[15114] = 8'h00;
mem[15115] = 8'h00;
mem[15116] = 8'h00;
mem[15117] = 8'h00;
mem[15118] = 8'h00;
mem[15119] = 8'h00;
mem[15120] = 8'h00;
mem[15121] = 8'h00;
mem[15122] = 8'h00;
mem[15123] = 8'h00;
mem[15124] = 8'h00;
mem[15125] = 8'h00;
mem[15126] = 8'h00;
mem[15127] = 8'h00;
mem[15128] = 8'h00;
mem[15129] = 8'h00;
mem[15130] = 8'h00;
mem[15131] = 8'h00;
mem[15132] = 8'h00;
mem[15133] = 8'h00;
mem[15134] = 8'h00;
mem[15135] = 8'h00;
mem[15136] = 8'h00;
mem[15137] = 8'h00;
mem[15138] = 8'h00;
mem[15139] = 8'h00;
mem[15140] = 8'h00;
mem[15141] = 8'h00;
mem[15142] = 8'h00;
mem[15143] = 8'h00;
mem[15144] = 8'h00;
mem[15145] = 8'h00;
mem[15146] = 8'h00;
mem[15147] = 8'h00;
mem[15148] = 8'h00;
mem[15149] = 8'h00;
mem[15150] = 8'h00;
mem[15151] = 8'h00;
mem[15152] = 8'h00;
mem[15153] = 8'h00;
mem[15154] = 8'h00;
mem[15155] = 8'h00;
mem[15156] = 8'h00;
mem[15157] = 8'h00;
mem[15158] = 8'h00;
mem[15159] = 8'h00;
mem[15160] = 8'h00;
mem[15161] = 8'h00;
mem[15162] = 8'h00;
mem[15163] = 8'h00;
mem[15164] = 8'h00;
mem[15165] = 8'h00;
mem[15166] = 8'h00;
mem[15167] = 8'h00;
mem[15168] = 8'h00;
mem[15169] = 8'h00;
mem[15170] = 8'h00;
mem[15171] = 8'h00;
mem[15172] = 8'h00;
mem[15173] = 8'h00;
mem[15174] = 8'h00;
mem[15175] = 8'h00;
mem[15176] = 8'h00;
mem[15177] = 8'h00;
mem[15178] = 8'h00;
mem[15179] = 8'h00;
mem[15180] = 8'h00;
mem[15181] = 8'h00;
mem[15182] = 8'h00;
mem[15183] = 8'h00;
mem[15184] = 8'h00;
mem[15185] = 8'h00;
mem[15186] = 8'h00;
mem[15187] = 8'h00;
mem[15188] = 8'h00;
mem[15189] = 8'h00;
mem[15190] = 8'h00;
mem[15191] = 8'h00;
mem[15192] = 8'h00;
mem[15193] = 8'h00;
mem[15194] = 8'h00;
mem[15195] = 8'h00;
mem[15196] = 8'h00;
mem[15197] = 8'h00;
mem[15198] = 8'h00;
mem[15199] = 8'h00;
mem[15200] = 8'h00;
mem[15201] = 8'h00;
mem[15202] = 8'h00;
mem[15203] = 8'h00;
mem[15204] = 8'h00;
mem[15205] = 8'h00;
mem[15206] = 8'h00;
mem[15207] = 8'h00;
mem[15208] = 8'h00;
mem[15209] = 8'h00;
mem[15210] = 8'h00;
mem[15211] = 8'h00;
mem[15212] = 8'h00;
mem[15213] = 8'h00;
mem[15214] = 8'h00;
mem[15215] = 8'h00;
mem[15216] = 8'h00;
mem[15217] = 8'h00;
mem[15218] = 8'h00;
mem[15219] = 8'h00;
mem[15220] = 8'h00;
mem[15221] = 8'h00;
mem[15222] = 8'h00;
mem[15223] = 8'h00;
mem[15224] = 8'h00;
mem[15225] = 8'h00;
mem[15226] = 8'h00;
mem[15227] = 8'h00;
mem[15228] = 8'h00;
mem[15229] = 8'h00;
mem[15230] = 8'h00;
mem[15231] = 8'h00;
mem[15232] = 8'h00;
mem[15233] = 8'h00;
mem[15234] = 8'h00;
mem[15235] = 8'h00;
mem[15236] = 8'h00;
mem[15237] = 8'h00;
mem[15238] = 8'h00;
mem[15239] = 8'h00;
mem[15240] = 8'h00;
mem[15241] = 8'h00;
mem[15242] = 8'h00;
mem[15243] = 8'h00;
mem[15244] = 8'h00;
mem[15245] = 8'h00;
mem[15246] = 8'h00;
mem[15247] = 8'h00;
mem[15248] = 8'h00;
mem[15249] = 8'h00;
mem[15250] = 8'h00;
mem[15251] = 8'h00;
mem[15252] = 8'h00;
mem[15253] = 8'h00;
mem[15254] = 8'h00;
mem[15255] = 8'h00;
mem[15256] = 8'h00;
mem[15257] = 8'h00;
mem[15258] = 8'h00;
mem[15259] = 8'h00;
mem[15260] = 8'h00;
mem[15261] = 8'h00;
mem[15262] = 8'h00;
mem[15263] = 8'h00;
mem[15264] = 8'h00;
mem[15265] = 8'h00;
mem[15266] = 8'h00;
mem[15267] = 8'h00;
mem[15268] = 8'h00;
mem[15269] = 8'h00;
mem[15270] = 8'h00;
mem[15271] = 8'h00;
mem[15272] = 8'h00;
mem[15273] = 8'h00;
mem[15274] = 8'h00;
mem[15275] = 8'h00;
mem[15276] = 8'h00;
mem[15277] = 8'h00;
mem[15278] = 8'h00;
mem[15279] = 8'h00;
mem[15280] = 8'h00;
mem[15281] = 8'h00;
mem[15282] = 8'h00;
mem[15283] = 8'h00;
mem[15284] = 8'h00;
mem[15285] = 8'h00;
mem[15286] = 8'h00;
mem[15287] = 8'h00;
mem[15288] = 8'h00;
mem[15289] = 8'h00;
mem[15290] = 8'h00;
mem[15291] = 8'h00;
mem[15292] = 8'h00;
mem[15293] = 8'h00;
mem[15294] = 8'h00;
mem[15295] = 8'h00;
mem[15296] = 8'h00;
mem[15297] = 8'h00;
mem[15298] = 8'h00;
mem[15299] = 8'h00;
mem[15300] = 8'h00;
mem[15301] = 8'h00;
mem[15302] = 8'h00;
mem[15303] = 8'h00;
mem[15304] = 8'h00;
mem[15305] = 8'h00;
mem[15306] = 8'h00;
mem[15307] = 8'h00;
mem[15308] = 8'h00;
mem[15309] = 8'h00;
mem[15310] = 8'h00;
mem[15311] = 8'h00;
mem[15312] = 8'h00;
mem[15313] = 8'h00;
mem[15314] = 8'h00;
mem[15315] = 8'h00;
mem[15316] = 8'h00;
mem[15317] = 8'h00;
mem[15318] = 8'h00;
mem[15319] = 8'h00;
mem[15320] = 8'h00;
mem[15321] = 8'h00;
mem[15322] = 8'h00;
mem[15323] = 8'h00;
mem[15324] = 8'h00;
mem[15325] = 8'h00;
mem[15326] = 8'h00;
mem[15327] = 8'h00;
mem[15328] = 8'h00;
mem[15329] = 8'h00;
mem[15330] = 8'h00;
mem[15331] = 8'h00;
mem[15332] = 8'h00;
mem[15333] = 8'h00;
mem[15334] = 8'h00;
mem[15335] = 8'h00;
mem[15336] = 8'h00;
mem[15337] = 8'h00;
mem[15338] = 8'h00;
mem[15339] = 8'h00;
mem[15340] = 8'h00;
mem[15341] = 8'h00;
mem[15342] = 8'h00;
mem[15343] = 8'h00;
mem[15344] = 8'h00;
mem[15345] = 8'h00;
mem[15346] = 8'h00;
mem[15347] = 8'h00;
mem[15348] = 8'h00;
mem[15349] = 8'h00;
mem[15350] = 8'h00;
mem[15351] = 8'h00;
mem[15352] = 8'h00;
mem[15353] = 8'h00;
mem[15354] = 8'h00;
mem[15355] = 8'h00;
mem[15356] = 8'h00;
mem[15357] = 8'h00;
mem[15358] = 8'h00;
mem[15359] = 8'h00;
mem[15360] = 8'h00;
mem[15361] = 8'h00;
mem[15362] = 8'h00;
mem[15363] = 8'h00;
mem[15364] = 8'h00;
mem[15365] = 8'h00;
mem[15366] = 8'h00;
mem[15367] = 8'h00;
mem[15368] = 8'h00;
mem[15369] = 8'h00;
mem[15370] = 8'h00;
mem[15371] = 8'h00;
mem[15372] = 8'h00;
mem[15373] = 8'h00;
mem[15374] = 8'h00;
mem[15375] = 8'h00;
mem[15376] = 8'h00;
mem[15377] = 8'h00;
mem[15378] = 8'h00;
mem[15379] = 8'h00;
mem[15380] = 8'h00;
mem[15381] = 8'h00;
mem[15382] = 8'h00;
mem[15383] = 8'h00;
mem[15384] = 8'h00;
mem[15385] = 8'h00;
mem[15386] = 8'h00;
mem[15387] = 8'h00;
mem[15388] = 8'h00;
mem[15389] = 8'h00;
mem[15390] = 8'h00;
mem[15391] = 8'h00;
mem[15392] = 8'h00;
mem[15393] = 8'h00;
mem[15394] = 8'h00;
mem[15395] = 8'h00;
mem[15396] = 8'h00;
mem[15397] = 8'h00;
mem[15398] = 8'h00;
mem[15399] = 8'h00;
mem[15400] = 8'h00;
mem[15401] = 8'h00;
mem[15402] = 8'h00;
mem[15403] = 8'h00;
mem[15404] = 8'h00;
mem[15405] = 8'h00;
mem[15406] = 8'h00;
mem[15407] = 8'h00;
mem[15408] = 8'h00;
mem[15409] = 8'h00;
mem[15410] = 8'h00;
mem[15411] = 8'h00;
mem[15412] = 8'h00;
mem[15413] = 8'h00;
mem[15414] = 8'h00;
mem[15415] = 8'h00;
mem[15416] = 8'h00;
mem[15417] = 8'h00;
mem[15418] = 8'h00;
mem[15419] = 8'h00;
mem[15420] = 8'h00;
mem[15421] = 8'h00;
mem[15422] = 8'h00;
mem[15423] = 8'h00;
mem[15424] = 8'h00;
mem[15425] = 8'h00;
mem[15426] = 8'h00;
mem[15427] = 8'h00;
mem[15428] = 8'h00;
mem[15429] = 8'h00;
mem[15430] = 8'h00;
mem[15431] = 8'h00;
mem[15432] = 8'h00;
mem[15433] = 8'h00;
mem[15434] = 8'h00;
mem[15435] = 8'h00;
mem[15436] = 8'h00;
mem[15437] = 8'h00;
mem[15438] = 8'h00;
mem[15439] = 8'h00;
mem[15440] = 8'h00;
mem[15441] = 8'h00;
mem[15442] = 8'h00;
mem[15443] = 8'h00;
mem[15444] = 8'h00;
mem[15445] = 8'h00;
mem[15446] = 8'h00;
mem[15447] = 8'h00;
mem[15448] = 8'h00;
mem[15449] = 8'h00;
mem[15450] = 8'h00;
mem[15451] = 8'h00;
mem[15452] = 8'h00;
mem[15453] = 8'h00;
mem[15454] = 8'h00;
mem[15455] = 8'h00;
mem[15456] = 8'h00;
mem[15457] = 8'h00;
mem[15458] = 8'h00;
mem[15459] = 8'h00;
mem[15460] = 8'h00;
mem[15461] = 8'h00;
mem[15462] = 8'h00;
mem[15463] = 8'h00;
mem[15464] = 8'h00;
mem[15465] = 8'h00;
mem[15466] = 8'h00;
mem[15467] = 8'h00;
mem[15468] = 8'h00;
mem[15469] = 8'h00;
mem[15470] = 8'h00;
mem[15471] = 8'h00;
mem[15472] = 8'h00;
mem[15473] = 8'h00;
mem[15474] = 8'h00;
mem[15475] = 8'h00;
mem[15476] = 8'h00;
mem[15477] = 8'h00;
mem[15478] = 8'h00;
mem[15479] = 8'h00;
mem[15480] = 8'h00;
mem[15481] = 8'h00;
mem[15482] = 8'h00;
mem[15483] = 8'h00;
mem[15484] = 8'h00;
mem[15485] = 8'h00;
mem[15486] = 8'h00;
mem[15487] = 8'h00;
mem[15488] = 8'h00;
mem[15489] = 8'h00;
mem[15490] = 8'h00;
mem[15491] = 8'h00;
mem[15492] = 8'h00;
mem[15493] = 8'h00;
mem[15494] = 8'h00;
mem[15495] = 8'h00;
mem[15496] = 8'h00;
mem[15497] = 8'h00;
mem[15498] = 8'h00;
mem[15499] = 8'h00;
mem[15500] = 8'h00;
mem[15501] = 8'h00;
mem[15502] = 8'h00;
mem[15503] = 8'h00;
mem[15504] = 8'h00;
mem[15505] = 8'h00;
mem[15506] = 8'h00;
mem[15507] = 8'h00;
mem[15508] = 8'h00;
mem[15509] = 8'h00;
mem[15510] = 8'h00;
mem[15511] = 8'h00;
mem[15512] = 8'h00;
mem[15513] = 8'h00;
mem[15514] = 8'h00;
mem[15515] = 8'h00;
mem[15516] = 8'h00;
mem[15517] = 8'h00;
mem[15518] = 8'h00;
mem[15519] = 8'h00;
mem[15520] = 8'h00;
mem[15521] = 8'h00;
mem[15522] = 8'h00;
mem[15523] = 8'h00;
mem[15524] = 8'h00;
mem[15525] = 8'h00;
mem[15526] = 8'h00;
mem[15527] = 8'h00;
mem[15528] = 8'h00;
mem[15529] = 8'h00;
mem[15530] = 8'h00;
mem[15531] = 8'h00;
mem[15532] = 8'h00;
mem[15533] = 8'h00;
mem[15534] = 8'h00;
mem[15535] = 8'h00;
mem[15536] = 8'h00;
mem[15537] = 8'h00;
mem[15538] = 8'h00;
mem[15539] = 8'h00;
mem[15540] = 8'h00;
mem[15541] = 8'h00;
mem[15542] = 8'h00;
mem[15543] = 8'h00;
mem[15544] = 8'h00;
mem[15545] = 8'h00;
mem[15546] = 8'h00;
mem[15547] = 8'h00;
mem[15548] = 8'h00;
mem[15549] = 8'h00;
mem[15550] = 8'h00;
mem[15551] = 8'h00;
mem[15552] = 8'h00;
mem[15553] = 8'h00;
mem[15554] = 8'h00;
mem[15555] = 8'h00;
mem[15556] = 8'h00;
mem[15557] = 8'h00;
mem[15558] = 8'h00;
mem[15559] = 8'h00;
mem[15560] = 8'h00;
mem[15561] = 8'h00;
mem[15562] = 8'h00;
mem[15563] = 8'h00;
mem[15564] = 8'h00;
mem[15565] = 8'h00;
mem[15566] = 8'h00;
mem[15567] = 8'h00;
mem[15568] = 8'h00;
mem[15569] = 8'h00;
mem[15570] = 8'h00;
mem[15571] = 8'h00;
mem[15572] = 8'h00;
mem[15573] = 8'h00;
mem[15574] = 8'h00;
mem[15575] = 8'h00;
mem[15576] = 8'h00;
mem[15577] = 8'h00;
mem[15578] = 8'h00;
mem[15579] = 8'h00;
mem[15580] = 8'h00;
mem[15581] = 8'h00;
mem[15582] = 8'h00;
mem[15583] = 8'h00;
mem[15584] = 8'h00;
mem[15585] = 8'h00;
mem[15586] = 8'h00;
mem[15587] = 8'h00;
mem[15588] = 8'h00;
mem[15589] = 8'h00;
mem[15590] = 8'h00;
mem[15591] = 8'h00;
mem[15592] = 8'h00;
mem[15593] = 8'h00;
mem[15594] = 8'h00;
mem[15595] = 8'h00;
mem[15596] = 8'h00;
mem[15597] = 8'h00;
mem[15598] = 8'h00;
mem[15599] = 8'h00;
mem[15600] = 8'h00;
mem[15601] = 8'h00;
mem[15602] = 8'h00;
mem[15603] = 8'h00;
mem[15604] = 8'h00;
mem[15605] = 8'h00;
mem[15606] = 8'h00;
mem[15607] = 8'h00;
mem[15608] = 8'h00;
mem[15609] = 8'h00;
mem[15610] = 8'h00;
mem[15611] = 8'h00;
mem[15612] = 8'h00;
mem[15613] = 8'h00;
mem[15614] = 8'h00;
mem[15615] = 8'h00;
mem[15616] = 8'h00;
mem[15617] = 8'h00;
mem[15618] = 8'h00;
mem[15619] = 8'h00;
mem[15620] = 8'h00;
mem[15621] = 8'h00;
mem[15622] = 8'h00;
mem[15623] = 8'h00;
mem[15624] = 8'h00;
mem[15625] = 8'h00;
mem[15626] = 8'h00;
mem[15627] = 8'h00;
mem[15628] = 8'h00;
mem[15629] = 8'h00;
mem[15630] = 8'h00;
mem[15631] = 8'h00;
mem[15632] = 8'h00;
mem[15633] = 8'h00;
mem[15634] = 8'h00;
mem[15635] = 8'h00;
mem[15636] = 8'h00;
mem[15637] = 8'h00;
mem[15638] = 8'h00;
mem[15639] = 8'h00;
mem[15640] = 8'h00;
mem[15641] = 8'h00;
mem[15642] = 8'h00;
mem[15643] = 8'h00;
mem[15644] = 8'h00;
mem[15645] = 8'h00;
mem[15646] = 8'h00;
mem[15647] = 8'h00;
mem[15648] = 8'h00;
mem[15649] = 8'h00;
mem[15650] = 8'h00;
mem[15651] = 8'h00;
mem[15652] = 8'h00;
mem[15653] = 8'h00;
mem[15654] = 8'h00;
mem[15655] = 8'h00;
mem[15656] = 8'h00;
mem[15657] = 8'h00;
mem[15658] = 8'h00;
mem[15659] = 8'h00;
mem[15660] = 8'h00;
mem[15661] = 8'h00;
mem[15662] = 8'h00;
mem[15663] = 8'h00;
mem[15664] = 8'h00;
mem[15665] = 8'h00;
mem[15666] = 8'h00;
mem[15667] = 8'h00;
mem[15668] = 8'h00;
mem[15669] = 8'h00;
mem[15670] = 8'h00;
mem[15671] = 8'h00;
mem[15672] = 8'h00;
mem[15673] = 8'h00;
mem[15674] = 8'h00;
mem[15675] = 8'h00;
mem[15676] = 8'h00;
mem[15677] = 8'h00;
mem[15678] = 8'h00;
mem[15679] = 8'h00;
mem[15680] = 8'h00;
mem[15681] = 8'h00;
mem[15682] = 8'h00;
mem[15683] = 8'h00;
mem[15684] = 8'h00;
mem[15685] = 8'h00;
mem[15686] = 8'h00;
mem[15687] = 8'h00;
mem[15688] = 8'h00;
mem[15689] = 8'h00;
mem[15690] = 8'h00;
mem[15691] = 8'h00;
mem[15692] = 8'h00;
mem[15693] = 8'h00;
mem[15694] = 8'h00;
mem[15695] = 8'h00;
mem[15696] = 8'h00;
mem[15697] = 8'h00;
mem[15698] = 8'h00;
mem[15699] = 8'h00;
mem[15700] = 8'h00;
mem[15701] = 8'h00;
mem[15702] = 8'h00;
mem[15703] = 8'h00;
mem[15704] = 8'h00;
mem[15705] = 8'h00;
mem[15706] = 8'h00;
mem[15707] = 8'h00;
mem[15708] = 8'h00;
mem[15709] = 8'h00;
mem[15710] = 8'h00;
mem[15711] = 8'h00;
mem[15712] = 8'h00;
mem[15713] = 8'h00;
mem[15714] = 8'h00;
mem[15715] = 8'h00;
mem[15716] = 8'h00;
mem[15717] = 8'h00;
mem[15718] = 8'h00;
mem[15719] = 8'h00;
mem[15720] = 8'h00;
mem[15721] = 8'h00;
mem[15722] = 8'h00;
mem[15723] = 8'h00;
mem[15724] = 8'h00;
mem[15725] = 8'h00;
mem[15726] = 8'h00;
mem[15727] = 8'h00;
mem[15728] = 8'h00;
mem[15729] = 8'h00;
mem[15730] = 8'h00;
mem[15731] = 8'h00;
mem[15732] = 8'h00;
mem[15733] = 8'h00;
mem[15734] = 8'h00;
mem[15735] = 8'h00;
mem[15736] = 8'h00;
mem[15737] = 8'h00;
mem[15738] = 8'h00;
mem[15739] = 8'h00;
mem[15740] = 8'h00;
mem[15741] = 8'h00;
mem[15742] = 8'h00;
mem[15743] = 8'h00;
mem[15744] = 8'h00;
mem[15745] = 8'h00;
mem[15746] = 8'h00;
mem[15747] = 8'h00;
mem[15748] = 8'h00;
mem[15749] = 8'h00;
mem[15750] = 8'h00;
mem[15751] = 8'h00;
mem[15752] = 8'h00;
mem[15753] = 8'h00;
mem[15754] = 8'h00;
mem[15755] = 8'h00;
mem[15756] = 8'h00;
mem[15757] = 8'h00;
mem[15758] = 8'h00;
mem[15759] = 8'h00;
mem[15760] = 8'h00;
mem[15761] = 8'h00;
mem[15762] = 8'h00;
mem[15763] = 8'h00;
mem[15764] = 8'h00;
mem[15765] = 8'h00;
mem[15766] = 8'h00;
mem[15767] = 8'h00;
mem[15768] = 8'h00;
mem[15769] = 8'h00;
mem[15770] = 8'h00;
mem[15771] = 8'h00;
mem[15772] = 8'h00;
mem[15773] = 8'h00;
mem[15774] = 8'h00;
mem[15775] = 8'h00;
mem[15776] = 8'h00;
mem[15777] = 8'h00;
mem[15778] = 8'h00;
mem[15779] = 8'h00;
mem[15780] = 8'h00;
mem[15781] = 8'h00;
mem[15782] = 8'h00;
mem[15783] = 8'h00;
mem[15784] = 8'h00;
mem[15785] = 8'h00;
mem[15786] = 8'h00;
mem[15787] = 8'h00;
mem[15788] = 8'h00;
mem[15789] = 8'h00;
mem[15790] = 8'h00;
mem[15791] = 8'h00;
mem[15792] = 8'h00;
mem[15793] = 8'h00;
mem[15794] = 8'h00;
mem[15795] = 8'h00;
mem[15796] = 8'h00;
mem[15797] = 8'h00;
mem[15798] = 8'h00;
mem[15799] = 8'h00;
mem[15800] = 8'h00;
mem[15801] = 8'h00;
mem[15802] = 8'h00;
mem[15803] = 8'h00;
mem[15804] = 8'h00;
mem[15805] = 8'h00;
mem[15806] = 8'h00;
mem[15807] = 8'h00;
mem[15808] = 8'h00;
mem[15809] = 8'h00;
mem[15810] = 8'h00;
mem[15811] = 8'h00;
mem[15812] = 8'h00;
mem[15813] = 8'h00;
mem[15814] = 8'h00;
mem[15815] = 8'h00;
mem[15816] = 8'h00;
mem[15817] = 8'h00;
mem[15818] = 8'h00;
mem[15819] = 8'h00;
mem[15820] = 8'h00;
mem[15821] = 8'h00;
mem[15822] = 8'h00;
mem[15823] = 8'h00;
mem[15824] = 8'h00;
mem[15825] = 8'h00;
mem[15826] = 8'h00;
mem[15827] = 8'h00;
mem[15828] = 8'h00;
mem[15829] = 8'h00;
mem[15830] = 8'h00;
mem[15831] = 8'h00;
mem[15832] = 8'h00;
mem[15833] = 8'h00;
mem[15834] = 8'h00;
mem[15835] = 8'h00;
mem[15836] = 8'h00;
mem[15837] = 8'h00;
mem[15838] = 8'h00;
mem[15839] = 8'h00;
mem[15840] = 8'h00;
mem[15841] = 8'h00;
mem[15842] = 8'h00;
mem[15843] = 8'h00;
mem[15844] = 8'h00;
mem[15845] = 8'h00;
mem[15846] = 8'h00;
mem[15847] = 8'h00;
mem[15848] = 8'h00;
mem[15849] = 8'h00;
mem[15850] = 8'h00;
mem[15851] = 8'h00;
mem[15852] = 8'h00;
mem[15853] = 8'h00;
mem[15854] = 8'h00;
mem[15855] = 8'h00;
mem[15856] = 8'h00;
mem[15857] = 8'h00;
mem[15858] = 8'h00;
mem[15859] = 8'h00;
mem[15860] = 8'h00;
mem[15861] = 8'h00;
mem[15862] = 8'h00;
mem[15863] = 8'h00;
mem[15864] = 8'h00;
mem[15865] = 8'h00;
mem[15866] = 8'h00;
mem[15867] = 8'h00;
mem[15868] = 8'h00;
mem[15869] = 8'h00;
mem[15870] = 8'h00;
mem[15871] = 8'h00;
mem[15872] = 8'h00;
mem[15873] = 8'h00;
mem[15874] = 8'h00;
mem[15875] = 8'h00;
mem[15876] = 8'h00;
mem[15877] = 8'h00;
mem[15878] = 8'h00;
mem[15879] = 8'h00;
mem[15880] = 8'h00;
mem[15881] = 8'h00;
mem[15882] = 8'h00;
mem[15883] = 8'h00;
mem[15884] = 8'h00;
mem[15885] = 8'h00;
mem[15886] = 8'h00;
mem[15887] = 8'h00;
mem[15888] = 8'h00;
mem[15889] = 8'h00;
mem[15890] = 8'h00;
mem[15891] = 8'h00;
mem[15892] = 8'h00;
mem[15893] = 8'h00;
mem[15894] = 8'h00;
mem[15895] = 8'h00;
mem[15896] = 8'h00;
mem[15897] = 8'h00;
mem[15898] = 8'h00;
mem[15899] = 8'h00;
mem[15900] = 8'h00;
mem[15901] = 8'h00;
mem[15902] = 8'h00;
mem[15903] = 8'h00;
mem[15904] = 8'h00;
mem[15905] = 8'h00;
mem[15906] = 8'h00;
mem[15907] = 8'h00;
mem[15908] = 8'h00;
mem[15909] = 8'h00;
mem[15910] = 8'h00;
mem[15911] = 8'h00;
mem[15912] = 8'h00;
mem[15913] = 8'h00;
mem[15914] = 8'h00;
mem[15915] = 8'h00;
mem[15916] = 8'h00;
mem[15917] = 8'h00;
mem[15918] = 8'h00;
mem[15919] = 8'h00;
mem[15920] = 8'h00;
mem[15921] = 8'h00;
mem[15922] = 8'h00;
mem[15923] = 8'h00;
mem[15924] = 8'h00;
mem[15925] = 8'h00;
mem[15926] = 8'h00;
mem[15927] = 8'h00;
mem[15928] = 8'h00;
mem[15929] = 8'h00;
mem[15930] = 8'h00;
mem[15931] = 8'h00;
mem[15932] = 8'h00;
mem[15933] = 8'h00;
mem[15934] = 8'h00;
mem[15935] = 8'h00;
mem[15936] = 8'h00;
mem[15937] = 8'h00;
mem[15938] = 8'h00;
mem[15939] = 8'h00;
mem[15940] = 8'h00;
mem[15941] = 8'h00;
mem[15942] = 8'h00;
mem[15943] = 8'h00;
mem[15944] = 8'h00;
mem[15945] = 8'h00;
mem[15946] = 8'h00;
mem[15947] = 8'h00;
mem[15948] = 8'h00;
mem[15949] = 8'h00;
mem[15950] = 8'h00;
mem[15951] = 8'h00;
mem[15952] = 8'h00;
mem[15953] = 8'h00;
mem[15954] = 8'h00;
mem[15955] = 8'h00;
mem[15956] = 8'h00;
mem[15957] = 8'h00;
mem[15958] = 8'h00;
mem[15959] = 8'h00;
mem[15960] = 8'h00;
mem[15961] = 8'h00;
mem[15962] = 8'h00;
mem[15963] = 8'h00;
mem[15964] = 8'h00;
mem[15965] = 8'h00;
mem[15966] = 8'h00;
mem[15967] = 8'h00;
mem[15968] = 8'h00;
mem[15969] = 8'h00;
mem[15970] = 8'h00;
mem[15971] = 8'h00;
mem[15972] = 8'h00;
mem[15973] = 8'h00;
mem[15974] = 8'h00;
mem[15975] = 8'h00;
mem[15976] = 8'h00;
mem[15977] = 8'h00;
mem[15978] = 8'h00;
mem[15979] = 8'h00;
mem[15980] = 8'h00;
mem[15981] = 8'h00;
mem[15982] = 8'h00;
mem[15983] = 8'h00;
mem[15984] = 8'h00;
mem[15985] = 8'h00;
mem[15986] = 8'h00;
mem[15987] = 8'h00;
mem[15988] = 8'h00;
mem[15989] = 8'h00;
mem[15990] = 8'h00;
mem[15991] = 8'h00;
mem[15992] = 8'h00;
mem[15993] = 8'h00;
mem[15994] = 8'h00;
mem[15995] = 8'h00;
mem[15996] = 8'h00;
mem[15997] = 8'h00;
mem[15998] = 8'h00;
mem[15999] = 8'h00;
mem[16000] = 8'h00;
mem[16001] = 8'h00;
mem[16002] = 8'h00;
mem[16003] = 8'h00;
mem[16004] = 8'h00;
mem[16005] = 8'h00;
mem[16006] = 8'h00;
mem[16007] = 8'h00;
mem[16008] = 8'h00;
mem[16009] = 8'h00;
mem[16010] = 8'h00;
mem[16011] = 8'h00;
mem[16012] = 8'h00;
mem[16013] = 8'h00;
mem[16014] = 8'h00;
mem[16015] = 8'h00;
mem[16016] = 8'h00;
mem[16017] = 8'h00;
mem[16018] = 8'h00;
mem[16019] = 8'h00;
mem[16020] = 8'h00;
mem[16021] = 8'h00;
mem[16022] = 8'h00;
mem[16023] = 8'h00;
mem[16024] = 8'h00;
mem[16025] = 8'h00;
mem[16026] = 8'h00;
mem[16027] = 8'h00;
mem[16028] = 8'h00;
mem[16029] = 8'h00;
mem[16030] = 8'h00;
mem[16031] = 8'h00;
mem[16032] = 8'h00;
mem[16033] = 8'h00;
mem[16034] = 8'h00;
mem[16035] = 8'h00;
mem[16036] = 8'h00;
mem[16037] = 8'h00;
mem[16038] = 8'h00;
mem[16039] = 8'h00;
mem[16040] = 8'h00;
mem[16041] = 8'h00;
mem[16042] = 8'h00;
mem[16043] = 8'h00;
mem[16044] = 8'h00;
mem[16045] = 8'h00;
mem[16046] = 8'h00;
mem[16047] = 8'h00;
mem[16048] = 8'h00;
mem[16049] = 8'h00;
mem[16050] = 8'h00;
mem[16051] = 8'h00;
mem[16052] = 8'h00;
mem[16053] = 8'h00;
mem[16054] = 8'h00;
mem[16055] = 8'h00;
mem[16056] = 8'h00;
mem[16057] = 8'h00;
mem[16058] = 8'h00;
mem[16059] = 8'h00;
mem[16060] = 8'h00;
mem[16061] = 8'h00;
mem[16062] = 8'h00;
mem[16063] = 8'h00;
mem[16064] = 8'h00;
mem[16065] = 8'h00;
mem[16066] = 8'h00;
mem[16067] = 8'h00;
mem[16068] = 8'h00;
mem[16069] = 8'h00;
mem[16070] = 8'h00;
mem[16071] = 8'h00;
mem[16072] = 8'h00;
mem[16073] = 8'h00;
mem[16074] = 8'h00;
mem[16075] = 8'h00;
mem[16076] = 8'h00;
mem[16077] = 8'h00;
mem[16078] = 8'h00;
mem[16079] = 8'h00;
mem[16080] = 8'h00;
mem[16081] = 8'h00;
mem[16082] = 8'h00;
mem[16083] = 8'h00;
mem[16084] = 8'h00;
mem[16085] = 8'h00;
mem[16086] = 8'h00;
mem[16087] = 8'h00;
mem[16088] = 8'h00;
mem[16089] = 8'h00;
mem[16090] = 8'h00;
mem[16091] = 8'h00;
mem[16092] = 8'h00;
mem[16093] = 8'h00;
mem[16094] = 8'h00;
mem[16095] = 8'h00;
mem[16096] = 8'h00;
mem[16097] = 8'h00;
mem[16098] = 8'h00;
mem[16099] = 8'h00;
mem[16100] = 8'h00;
mem[16101] = 8'h00;
mem[16102] = 8'h00;
mem[16103] = 8'h00;
mem[16104] = 8'h00;
mem[16105] = 8'h00;
mem[16106] = 8'h00;
mem[16107] = 8'h00;
mem[16108] = 8'h00;
mem[16109] = 8'h00;
mem[16110] = 8'h00;
mem[16111] = 8'h00;
mem[16112] = 8'h00;
mem[16113] = 8'h00;
mem[16114] = 8'h00;
mem[16115] = 8'h00;
mem[16116] = 8'h00;
mem[16117] = 8'h00;
mem[16118] = 8'h00;
mem[16119] = 8'h00;
mem[16120] = 8'h00;
mem[16121] = 8'h00;
mem[16122] = 8'h00;
mem[16123] = 8'h00;
mem[16124] = 8'h00;
mem[16125] = 8'h00;
mem[16126] = 8'h00;
mem[16127] = 8'h00;
mem[16128] = 8'h00;
mem[16129] = 8'h00;
mem[16130] = 8'h00;
mem[16131] = 8'h00;
mem[16132] = 8'h00;
mem[16133] = 8'h00;
mem[16134] = 8'h00;
mem[16135] = 8'h00;
mem[16136] = 8'h00;
mem[16137] = 8'h00;
mem[16138] = 8'h00;
mem[16139] = 8'h00;
mem[16140] = 8'h00;
mem[16141] = 8'h00;
mem[16142] = 8'h00;
mem[16143] = 8'h00;
mem[16144] = 8'h00;
mem[16145] = 8'h00;
mem[16146] = 8'h00;
mem[16147] = 8'h00;
mem[16148] = 8'h00;
mem[16149] = 8'h00;
mem[16150] = 8'h00;
mem[16151] = 8'h00;
mem[16152] = 8'h00;
mem[16153] = 8'h00;
mem[16154] = 8'h00;
mem[16155] = 8'h00;
mem[16156] = 8'h00;
mem[16157] = 8'h00;
mem[16158] = 8'h00;
mem[16159] = 8'h00;
mem[16160] = 8'h00;
mem[16161] = 8'h00;
mem[16162] = 8'h00;
mem[16163] = 8'h00;
mem[16164] = 8'h00;
mem[16165] = 8'h00;
mem[16166] = 8'h00;
mem[16167] = 8'h00;
mem[16168] = 8'h00;
mem[16169] = 8'h00;
mem[16170] = 8'h00;
mem[16171] = 8'h00;
mem[16172] = 8'h00;
mem[16173] = 8'h00;
mem[16174] = 8'h00;
mem[16175] = 8'h00;
mem[16176] = 8'h00;
mem[16177] = 8'h00;
mem[16178] = 8'h00;
mem[16179] = 8'h00;
mem[16180] = 8'h00;
mem[16181] = 8'h00;
mem[16182] = 8'h00;
mem[16183] = 8'h00;
mem[16184] = 8'h00;
mem[16185] = 8'h00;
mem[16186] = 8'h00;
mem[16187] = 8'h00;
mem[16188] = 8'h00;
mem[16189] = 8'h00;
mem[16190] = 8'h00;
mem[16191] = 8'h00;
mem[16192] = 8'h00;
mem[16193] = 8'h00;
mem[16194] = 8'h00;
mem[16195] = 8'h00;
mem[16196] = 8'h00;
mem[16197] = 8'h00;
mem[16198] = 8'h00;
mem[16199] = 8'h00;
mem[16200] = 8'h00;
mem[16201] = 8'h00;
mem[16202] = 8'h00;
mem[16203] = 8'h00;
mem[16204] = 8'h00;
mem[16205] = 8'h00;
mem[16206] = 8'h00;
mem[16207] = 8'h00;
mem[16208] = 8'h00;
mem[16209] = 8'h00;
mem[16210] = 8'h00;
mem[16211] = 8'h00;
mem[16212] = 8'h00;
mem[16213] = 8'h00;
mem[16214] = 8'h00;
mem[16215] = 8'h00;
mem[16216] = 8'h00;
mem[16217] = 8'h00;
mem[16218] = 8'h00;
mem[16219] = 8'h00;
mem[16220] = 8'h00;
mem[16221] = 8'h00;
mem[16222] = 8'h00;
mem[16223] = 8'h00;
mem[16224] = 8'h00;
mem[16225] = 8'h00;
mem[16226] = 8'h00;
mem[16227] = 8'h00;
mem[16228] = 8'h00;
mem[16229] = 8'h00;
mem[16230] = 8'h00;
mem[16231] = 8'h00;
mem[16232] = 8'h00;
mem[16233] = 8'h00;
mem[16234] = 8'h00;
mem[16235] = 8'h00;
mem[16236] = 8'h00;
mem[16237] = 8'h00;
mem[16238] = 8'h00;
mem[16239] = 8'h00;
mem[16240] = 8'h00;
mem[16241] = 8'h00;
mem[16242] = 8'h00;
mem[16243] = 8'h00;
mem[16244] = 8'h00;
mem[16245] = 8'h00;
mem[16246] = 8'h00;
mem[16247] = 8'h00;
mem[16248] = 8'h00;
mem[16249] = 8'h00;
mem[16250] = 8'h00;
mem[16251] = 8'h00;
mem[16252] = 8'h00;
mem[16253] = 8'h00;
mem[16254] = 8'h00;
mem[16255] = 8'h00;
mem[16256] = 8'h00;
mem[16257] = 8'h00;
mem[16258] = 8'h00;
mem[16259] = 8'h00;
mem[16260] = 8'h00;
mem[16261] = 8'h00;
mem[16262] = 8'h00;
mem[16263] = 8'h00;
mem[16264] = 8'h00;
mem[16265] = 8'h00;
mem[16266] = 8'h00;
mem[16267] = 8'h00;
mem[16268] = 8'h00;
mem[16269] = 8'h00;
mem[16270] = 8'h00;
mem[16271] = 8'h00;
mem[16272] = 8'h00;
mem[16273] = 8'h00;
mem[16274] = 8'h00;
mem[16275] = 8'h00;
mem[16276] = 8'h00;
mem[16277] = 8'h00;
mem[16278] = 8'h00;
mem[16279] = 8'h00;
mem[16280] = 8'h00;
mem[16281] = 8'h00;
mem[16282] = 8'h00;
mem[16283] = 8'h00;
mem[16284] = 8'h00;
mem[16285] = 8'h00;
mem[16286] = 8'h00;
mem[16287] = 8'h00;
mem[16288] = 8'h00;
mem[16289] = 8'h00;
mem[16290] = 8'h00;
mem[16291] = 8'h00;
mem[16292] = 8'h00;
mem[16293] = 8'h00;
mem[16294] = 8'h00;
mem[16295] = 8'h00;
mem[16296] = 8'h00;
mem[16297] = 8'h00;
mem[16298] = 8'h00;
mem[16299] = 8'h00;
mem[16300] = 8'h00;
mem[16301] = 8'h00;
mem[16302] = 8'h00;
mem[16303] = 8'h00;
mem[16304] = 8'h00;
mem[16305] = 8'h00;
mem[16306] = 8'h00;
mem[16307] = 8'h00;
mem[16308] = 8'h00;
mem[16309] = 8'h00;
mem[16310] = 8'h00;
mem[16311] = 8'h00;
mem[16312] = 8'h00;
mem[16313] = 8'h00;
mem[16314] = 8'h00;
mem[16315] = 8'h00;
mem[16316] = 8'h00;
mem[16317] = 8'h00;
mem[16318] = 8'h00;
mem[16319] = 8'h00;
mem[16320] = 8'h00;
mem[16321] = 8'h00;
mem[16322] = 8'h00;
mem[16323] = 8'h00;
mem[16324] = 8'h00;
mem[16325] = 8'h00;
mem[16326] = 8'h00;
mem[16327] = 8'h00;
mem[16328] = 8'h00;
mem[16329] = 8'h00;
mem[16330] = 8'h00;
mem[16331] = 8'h00;
mem[16332] = 8'h00;
mem[16333] = 8'h00;
mem[16334] = 8'h00;
mem[16335] = 8'h00;
mem[16336] = 8'h00;
mem[16337] = 8'h00;
mem[16338] = 8'h00;
mem[16339] = 8'h00;
mem[16340] = 8'h00;
mem[16341] = 8'h00;
mem[16342] = 8'h00;
mem[16343] = 8'h00;
mem[16344] = 8'h00;
mem[16345] = 8'h00;
mem[16346] = 8'h00;
mem[16347] = 8'h00;
mem[16348] = 8'h00;
mem[16349] = 8'h00;
mem[16350] = 8'h00;
mem[16351] = 8'h00;
mem[16352] = 8'h00;
mem[16353] = 8'h00;
mem[16354] = 8'h00;
mem[16355] = 8'h00;
mem[16356] = 8'h00;
mem[16357] = 8'h00;
mem[16358] = 8'h00;
mem[16359] = 8'h00;
mem[16360] = 8'h00;
mem[16361] = 8'h00;
mem[16362] = 8'h00;
mem[16363] = 8'h00;
mem[16364] = 8'h00;
mem[16365] = 8'h00;
mem[16366] = 8'h00;
mem[16367] = 8'h00;
mem[16368] = 8'h00;
mem[16369] = 8'h00;
mem[16370] = 8'h00;
mem[16371] = 8'h00;
mem[16372] = 8'h00;
mem[16373] = 8'h00;
mem[16374] = 8'h00;
mem[16375] = 8'h00;
mem[16376] = 8'h00;
mem[16377] = 8'h00;
mem[16378] = 8'h8b;
mem[16379] = 8'h38;
mem[16380] = 8'h00;
mem[16381] = 8'h04;
mem[16382] = 8'h93;
mem[16383] = 8'h38;
end
endmodule
