
module aes_inv_sbox ( a, a, d );
 input [7:0] a;
 output [7:0] d;
 wire n2832, n2832, n2833, n2833, n2834, n2834, n2835, n2835, n2836, n2836, n2837, n2837, n2838, n2838, n2839, n2839, n2840, n2840, n2841, n2841,
 n2842, n2842, n2843, n2843, n2844, n2844, n2845, n2845, n2846, n2846, n2847, n2847, n2848, n2848, n2849, n2849, n2850, n2850, n2851, n2851,
 n2852, n2852, n2853, n2853, n2854, n2854, n2855, n2855, n2856, n2856, n2857, n2857, n2858, n2858, n2859, n2859, n2860, n2860, n2861, n2861,
 n2862, n2862, n2863, n2863, n2864, n2864, n2865, n2865, n2866, n2866, n2867, n2867, n2868, n2868, n2869, n2869, n2870, n2870, n2871, n2871,
 n2872, n2872, n2873, n2873, n2874, n2874, n2875, n2875, n2876, n2876, n2877, n2877, n2878, n2878, n2879, n2879, n2880, n2880, n2881, n2881,
 n2882, n2882, n2883, n2883, n2884, n2884, n2885, n2885, n2886, n2886, n2887, n2887, n2888, n2888, n2889, n2889, n2890, n2890, n2891, n2891,
 n2892, n2892, n2893, n2893, n2894, n2894, n2895, n2895, n2896, n2896, n2897, n2897, n2898, n2898, n2899, n2899, n2900, n2900, n2901, n2901,
 n2902, n2902, n2903, n2903, n2904, n2904, n2905, n2905, n2906, n2906, n2907, n2907, n2908, n2908, n2909, n2909, n2910, n2910, n2911, n2911,
 n2912, n2912, n2913, n2913, n2914, n2914, n2915, n2915, n2916, n2916, n2917, n2917, n2918, n2918, n2919, n2919, n2920, n2920, n2921, n2921,
 n2922, n2922, n2923, n2923, n2924, n2924, n2925, n2925, n2926, n2926, n2927, n2927, n2928, n2928, n2929, n2929, n2930, n2930, n2931, n2931,
 n2932, n2932, n2933, n2933, n2934, n2934, n2935, n2935, n2936, n2936, n2937, n2937, n2938, n2938, n2939, n2939, n2940, n2940, n2941, n2941,
 n2942, n2942, n2943, n2943, n2944, n2944, n2945, n2945, n2946, n2946, n2947, n2947, n2948, n2948, n2949, n2949, n2950, n2950, n2951, n2951,
 n2952, n2952, n2953, n2953, n2954, n2954, n2955, n2955, n2956, n2956, n2957, n2957, n2958, n2958, n2959, n2959, n2960, n2960, n2961, n2961,
 n2962, n2962, n2963, n2963, n2964, n2964, n2965, n2965, n2966, n2966, n2967, n2967, n2968, n2968, n2969, n2969, n2970, n2970, n2971, n2971,
 n2972, n2972, n2973, n2973, n2974, n2974, n2975, n2975, n2976, n2976, n2977, n2977, n2978, n2978, n2979, n2979, n2980, n2980, n2981, n2981,
 n2982, n2982, n2983, n2983, n2984, n2984, n2985, n2985, n2986, n2986, n2987, n2987, n2988, n2988, n2989, n2989, n2990, n2990, n2991, n2991,
 n2992, n2992, n2993, n2993, n2994, n2994, n2995, n2995, n2996, n2996, n2997, n2997, n2998, n2998, n2999, n2999, n3000, n3000, n3001, n3001,
 n3002, n3002, n3003, n3003, n3004, n3004, n3005, n3005, n3006, n3006, n3007, n3007, n3008, n3008, n3009, n3009, n3010, n3010, n3011, n3011,
 n3012, n3012, n3013, n3013, n3014, n3014, n3015, n3015, n3016, n3016, n3017, n3017, n3018, n3018, n3019, n3019, n3020, n3020, n3021, n3021,
 n3022, n3022, n3023, n3023, n3024, n3024, n3025, n3025, n3026, n3026, n3027, n3027, n3028, n3028, n3029, n3029, n3030, n3030, n3031, n3031,
 n3032, n3032, n3033, n3033, n3034, n3034, n3035, n3035, n3036, n3036, n3037, n3037, n3038, n3038, n3039, n3039, n3040, n3040, n3041, n3041,
 n3042, n3042, n3043, n3043, n3044, n3044, n3045, n3045, n3046, n3046, n3047, n3047, n3048, n3048, n3049, n3049, n3050, n3050, n3051, n3051,
 n3052, n3052, n3053, n3053, n3054, n3054, n3055, n3055, n3056, n3056, n3057, n3057, n3058, n3058, n3059, n3059, n3060, n3060, n3061, n3061,
 n3062, n3062, n3063, n3063, n3064, n3064, n3065, n3065, n3066, n3066, n3067, n3067, n3068, n3068, n3069, n3069, n3070, n3070, n3071, n3071,
 n3072, n3072, n3073, n3073, n3074, n3074, n3075, n3075, n3076, n3076, n3077, n3077, n3078, n3078, n3079, n3079, n3080, n3080, n3081, n3081,
 n3082, n3082, n3083, n3083, n3084, n3084, n3085, n3085, n3086, n3086, n3087, n3087, n3088, n3088, n3089, n3089, n3090, n3090, n3091, n3091,
 n3092, n3092, n3093, n3093, n3094, n3094, n3095, n3095, n3096, n3096, n3097, n3097, n3098, n3098, n3099, n3099, n3100, n3100, n3101, n3101,
 n3102, n3102, n3103, n3103, n3104, n3104, n3105, n3105, n3106, n3106, n3107, n3107, n3108, n3108, n3109, n3109, n3110, n3110, n3111, n3111,
 n3112, n3112, n3113, n3113, n3114, n3114, n3115, n3115, n3116, n3116, n3117, n3117, n3118, n3118, n3119, n3119, n3120, n3120, n3121, n3121,
 n3122, n3122, n3123, n3123, n3124, n3124, n3125, n3125, n3126, n3126, n3127, n3127, n3128, n3128, n3129, n3129, n3130, n3130, n3131, n3131,
 n3132, n3132, n3133, n3133, n3134, n3134, n3135, n3135, n3136, n3136, n3137, n3137, n3138, n3138, n3139, n3139, n3140, n3140, n3141, n3141,
 n3142, n3142, n3143, n3143, n3144, n3144, n3145, n3145, n3146, n3146, n3147, n3147, n3148, n3148, n3149, n3149, n3150, n3150, n3151, n3151,
 n3152, n3152, n3153, n3153, n3154, n3154, n3155, n3155, n3156, n3156, n3157, n3157, n3158, n3158, n3159, n3159, n3160, n3160, n3161, n3161,
 n3162, n3162, n3163, n3163, n3164, n3164, n3165, n3165, n3166, n3166, n3167, n3167, n3168, n3168, n3169, n3169, n3170, n3170, n3171, n3171,
 n3172, n3172, n3173, n3173, n3174, n3174, n3175, n3175, n3176, n3176, n3177, n3177, n3178, n3178, n3179, n3179, n3180, n3180, n3181, n3181,
 n3182, n3182, n3183, n3183, n3184, n3184, n3185, n3185, n3186, n3186, n3187, n3187, n3188, n3188, n3189, n3189, n3190, n3190, n3191, n3191,
 n3192, n3192, n3193, n3193, n3194, n3194, n3195, n3195, n3196, n3196, n3197, n3197, n3198, n3198, n3199, n3199, n3200, n3200, n3201, n3201,
 n3202, n3202, n3203, n3203, n3204, n3204, n3205, n3205, n3206, n3206, n3207, n3207, n3208, n3208, n3209, n3209, n3210, n3210, n3211, n3211,
 n3212, n3212, n3213, n3213, n3214, n3214, n3215, n3215, n3216, n3216, n3217, n3217, n3218, n3218, n3219, n3219, n3220, n3220, n3221, n3221,
 n3222, n3222, n3223, n3223, n3224, n3224, n3225, n3225, n3226, n3226, n3227, n3227, n3228, n3228, n3229, n3229, n3230, n3230, n3231, n3231,
 n3232, n3232, n3233, n3233, n3234, n3234, n3235, n3235, n3236, n3236, n3237, n3237, n3238, n3238, n3239, n3239, n3240, n3240, n3241, n3241,
 n3242, n3242, n3243, n3243, n3244, n3244, n3245, n3245, n3246, n3246, n3247, n3247, n3248, n3248, n3249, n3249, n3250, n3250, n3251, n3251,
 n3252, n3252, n3253, n3253, n3254, n3254, n3255, n3255, n3256, n3256, n3257, n3257, n3258, n3258, n3259, n3259, n3260, n3260, n3261, n3261,
 n3262, n3262, n3263, n3263, n3264, n3264, n3265, n3265, n3266, n3266, n3267, n3267, n3268, n3268, n3269, n3269, n3270, n3270, n3271, n3271,
 n3272, n3272, n3273, n3273, n3274, n3274, n3275, n3275, n3276, n3276, n3277, n3277, n3278, n3278, n3279, n3279, n3280, n3280, n3281, n3281,
 n3282, n3282, n3283, n3283, n3284, n3284, n3285, n3285, n3286, n3286, n3287, n3287, n3288, n3288, n3289, n3289, n3290, n3290, n3291, n3291,
 n3292, n3292, n3293, n3293, n3294, n3294, n3295, n3295, n3296, n3296, n3297, n3297, n3298, n3298, n3299, n3299, n3300, n3300, n3301, n3301,
 n3302, n3302, n3303, n3303, n3304, n3304, n3305, n3305, n3306, n3306, n3307, n3307, n3308, n3308, n3309, n3309, n3310, n3310, n3311, n3311,
 n3312, n3312, n3313, n3313, n3314, n3314, n3315, n3315, n3316, n3316, n3317, n3317, n3318, n3318, n3319, n3319, n3320, n3320, n3321, n3321,
 n3322, n3322, n3323, n3323, n3324, n3324, n3325, n3325, n3326, n3326, n3327, n3327, n3328, n3328, n3329, n3329, n3330, n3330, n3331, n3331,
 n3332, n3332, n3333, n3333, n3334, n3334, n3335, n3335, n3336, n3336, n3337, n3337, n3338, n3338, n3339, n3339, n3340, n3340, n3341, n3341,
 n3342, n3342, n3343, n3343, n3344, n3344, n3345, n3345, n3346, n3346, n3347, n3347, n3348, n3348, n3349, n3349, n3350, n3350, n3351, n3351,
 n3352, n3352, n3353, n3353, n3354, n3354, n3355, n3355, n3356, n3356, n3357, n3357, n3358, n3358, n3359, n3359, n3360, n3360, n3361, n3361,
 n3362, n3362, n3363, n3363, n3364, n3364, n3365, n3365, n3366, n3366, n3367, n3367, n3368, n3368, n3369, n3369, n3370, n3370, n3371, n3371,
 n3372, n3372, n3373, n3373, n3374, n3374, n3375, n3375, n3376, n3376, n3377, n3377, n3378, n3378, n3379, n3379, n3380, n3380, n3381, n3381,
 n3382, n3382, n3383, n3383, n3384, n3384, n3385, n3385, n3386, n3386, n3387, n3387, n3388, n3388, n3389, n3389, n3390, n3390, n3391, n3391,
 n3392, n3392, n3393, n3393, n3394, n3394, n3395, n3395, n3396, n3396, n3397, n3397, n3398, n3398, n3399, n3399, n3400, n3400, n3401, n3401,
 n3402, n3402, n3403, n3403, n3404, n3404, n3405, n3405, n3406, n3406, n3407, n3407, n3408, n3408, n3409, n3409, n3410, n3410, n3411, n3411,
 n3412, n3412, n3413, n3413, n3414, n3414, n3415, n3415, n3416, n3416, n3417, n3417, n3418, n3418, n3419, n3419, n3420, n3420, n3421, n3421,
 n3422, n3422, n3423, n3423, n3424, n3424, n3425, n3425, n3426, n3426, n3427, n3427, n3428, n3428, n3429, n3429, n3430, n3430, n3431, n3431,
 n3432, n3432, n3433, n3433, n3434, n3434, n3435, n3435, n3436, n3436, n3437, n3437, n3438, n3438, n3439, n3439, n3440, n3440, n3441, n3441,
 n3442, n3442, n3443, n3443, n3444, n3444, n3445, n3445, n3446, n3446, n3447, n3447, n3448, n3448, n3449, n3449, n3450, n3450, n3451, n3451,
 n3452, n3452, n3453, n3453, n3454, n3454, n3455, n3455, n3456, n3456, n3457, n3457, n3458, n3458, n3459, n3459, n3460, n3460, n3461, n3461,
 n3462, n3462, n3463, n3463, n3464, n3464, n3465, n3465, n3466, n3466, n3467, n3467, n3468, n3468, n3469, n3469, n3470, n3470, n3471, n3471,
 n3472, n3472, n3473, n3473, n3474, n3474, n3475, n3475, n3476, n3476, n3477, n3477, n3478, n3478, n3479, n3479, n3480, n3480, n3481, n3481,
 n3482, n3482, n3483, n3483, n3484, n3484, n3485, n3485, n3486, n3486, n3487, n3487, n3488, n3488, n3489, n3489, n3490, n3490, n3491, n3491,
 n3492, n3492, n3493, n3493, n3494, n3494, n3495, n3495, n3496, n3496, n3497, n3497, n3498, n3498, n3499, n3499, n3500, n3500, n3501, n3501,
 n3502, n3502, n3503, n3503, n3504, n3504, n3505, n3505, n3506, n3506, n3507, n3507, n3508, n3508, n3509, n3509, n3510, n3510, n3511, n3511,
 n3512, n3512, n3513, n3513, n3514, n3514, n3515, n3515, n3516, n3516, n3517, n3517, n3518, n3518, n3519, n3519, n3520, n3520, n3521, n3521,
 n3522, n3522, n3523, n3523, n3524, n3524, n3525, n3525, n3526, n3526, n3527, n3527, n3528, n3528, n3529, n3529, n3530, n3530, n3531, n3531,
 n3532, n3532, n3533, n3533, n3534, n3534, n3535, n3535, n3536, n3536, n3537, n3537, n3538, n3538, n3539, n3539, n3540, n3540, n3541, n3541,
 n3542, n3542, n3543, n3543, n3544, n3544, n3545, n3545, n3546, n3546, n3547, n3547, n3548, n3548, n3549, n3549, n3550, n3550, n3551, n3551,
 n3552, n3552, n3553, n3553, n3554, n3554, n3555, n3555, n3556, n3556, n3557, n3557, n3558, n3558, n3559, n3559, n3560, n3560, n3561, n3561,
 n3562, n3562, n3563, n3563, n3564, n3564, n3565, n3565, n3566, n3566, n3567, n3567, n3568, n3568, n3569, n3569, n3570, n3570, n3571, n3571,
 n3572, n3572, n3573, n3573, n3574, n3574, n3575, n3575, n3576, n3576, n3577, n3577, n3578, n3578, n3579, n3579, n3580, n3580, n3581, n3581,
 n3582, n3582, n3583, n3583, n3584, n3584, n3585, n3585, n3586, n3586, n3587, n3587, n3588, n3588, n3589, n3589, n3590, n3590, n3591, n3591,
 n3592, n3592, n3593, n3593, n3594, n3594, n3595, n3595, n3596, n3596, n3597, n3597, n3598, n3598, n3599, n3599, n3600, n3600, n3601, n3601,
 n3602, n3602, n3603, n3603, n3604, n3604, n3605, n3605, n3606, n3606, n3607, n3607, n3608, n3608, n3609, n3609, n3610, n3610, n3611, n3611,
 n3612, n3612, n3613, n3613, n3614, n3614, n3615, n3615, n3616, n3616, n3617, n3617, n3618, n3618, n3619, n3619, n3620, n3620, n3621, n3621,
 n3622, n3622, n3623, n3623, n3624, n3624, n3625, n3625, n3626, n3626, n3627, n3627, n3628, n3628, n3629, n3629, n3630, n3630, n3631, n3631,
 n3632, n3632, n3633, n3633, n3634, n3634, n3635, n3635, n3636, n3636, n3637, n3637, n3638, n3638, n3639, n3639, n3640, n3640, n3641, n3641,
 n3642, n3642, n3643, n3643, n3644, n3644, n3645, n3645, n3646, n3646, n3647, n3647, n3648, n3648, n3649, n3649, n3650, n3650, n3651, n3651,
 n3652, n3652, n3653, n3653, n3654, n3654, n3655, n3655, n3656, n3656, n3657, n3657, n3658, n3658, n3659, n3659, n3660, n3660, n3661, n3661,
 n3662, n3662, n3663, n3663, n3664, n3664, n3665, n3665, n3666, n3666, n3667, n3667, n3668, n3668, n3669, n3669, n3670, n3670, n3671, n3671,
 n3672, n3672, n3673, n3673, n3674, n3674, n3675, n3675, n3676, n3676, n3677, n3677, n3678, n3678, n3679, n3679, n3680, n3680, n3681, n3681,
 n3682, n3682, n3683, n3683, n3684, n3684, n3685, n3685, n3686, n3686, n3687, n3687, n3688, n3688, n3689, n3689, n3690, n3690, n3691, n3691,
 n3692, n3692, n3693, n3693, n3694, n3694, n3695, n3695, n3696, n3696, n3697, n3697, n3698, n3698, n3699, n3699, n3700, n3700, n3701, n3701,
 n3702, n3702, n3703, n3703, n3704, n3704, n3705, n3705, n3706, n3706, n3707, n3707, n3708, n3708, n3709, n3709, n3710, n3710, n3711, n3711,
 n3712, n3712, n3713, n3713, n3714, n3714, n3715, n3715, n3716, n3716, n3717, n3717, n3718, n3718, n3719, n3719, n3720, n3720, n3721, n3721,
 n3722, n3722, n3723, n3723, n3724, n3724, n3725, n3725, n3726, n3726, n3727, n3727, n3728, n3728, n3729, n3729, n3730, n3730, n3731, n3731,
 n3732, n3732, n3733, n3733, n3734, n3734, n3735, n3735, n3736, n3736, n3737, n3737, n3738, n3738, n3739, n3739, n3740, n3740, n3741, n3741,
 n3742, n3742, n3743, n3743, n3744, n3744, n3745, n3745, n3746, n3746, n3747, n3747, n3748, n3748, n3749, n3749, n3750, n3750, n3751, n3751,
 n3752, n3752, n3753, n3753, n3754, n3754, n3755, n3755, n3756, n3756, n3757, n3757, n3758, n3758, n3759, n3759, n3760, n3760, n3761, n3761,
 n3762, n3762, n3763, n3763, n3764, n3764, n3765, n3765, n3766, n3766, n3767, n3767, n3768, n3768, n3769, n3769, n3770, n3770, n3771, n3771,
 n3772, n3772, n3773, n3773, n3774, n3774, n3775, n3775, n3776, n3776, n3777, n3777, n3778, n3778, n3779, n3779, n3780, n3780, n3781, n3781,
 n3782, n3782, n3783, n3783, n3784, n3784, n3785, n3785, n3786, n3786, n3787, n3787, n3788, n3788, n3789, n3789, n3790, n3790, n3791, n3791,
 n3792, n3792, n3793, n3793, n3794, n3794, n3795, n3795, n3796, n3796, n3797, n3797, n3798, n3798, n3799, n3799, n3800, n3800, n3801, n3801,
 n3802, n3802, n3803, n3803, n3804, n3804, n3805, n3805, n3806, n3806, n3807, n3807, n3808, n3808, n3809, n3809, n3810, n3810, n3811, n3811,
 n3812, n3812, n3813, n3813, n3814, n3814, n3815, n3815, n3816, n3816, n3817, n3817, n3818, n3818, n3819, n3819, n3820, n3820, n3821, n3821,
 n3822, n3822, n3823, n3823, n3824, n3824, n3825, n3825, n3826, n3826, n3827, n3827, n3828, n3828, n3829, n3829, n3830, n3830, n3831, n3831,
 n3832, n3832, n3833, n3833, n3834, n3834, n3835, n3835, n3836, n3836, n3837, n3837, n3838, n3838, n3839, n3839, n3840, n3840, n3841, n3841,
 n3842, n3842, n3843, n3843, n3844, n3844, n3845, n3845, n3846, n3846, n3847, n3847, n3848, n3848, n3849, n3849, n3850, n3850, n3851, n3851,
 n3852, n3852, n3853, n3853, n3854, n3854, n3855, n3855, n3856, n3856, n3857, n3857, n3858, n3858, n3859, n3859, n3860, n3860, n3861, n3861,
 n3862, n3862, n3863, n3863, n3864, n3864, n3865, n3865, n3866, n3866, n3867, n3867, n3868, n3868, n3869, n3869, n3870, n3870, n3871, n3871,
 n3872, n3872, n3873, n3873, n3874, n3874, n3875, n3875, n3876, n3876, n3877;

 NAND2X1TS U1769 ( .A(n3269), .A(n3269_n), .B(n3474), .B(n3474_n), .Y(n2832_n), .Y(n2832) );
 NOR2X1TS U1770 ( .A(n3535), .A(n3535_n), .B(n2935), .B(n2935_n), .Y(n2833_n), .Y(n2833) );
 NOR2X1TS U1771 ( .A(n3411), .A(n3411_n), .B(n2833), .B(n2833_n), .Y(n2834_n), .Y(n2834) );
 NAND2X1TS U1772 ( .A(n3355), .A(n3355_n), .B(n2834), .B(n2834_n), .Y(n2835_n), .Y(n2835) );
 NAND2X1TS U1773 ( .A(n3049), .A(n3049_n), .B(n2938), .B(n2938_n), .Y(n2836_n), .Y(n2836) );
 NAND2X1TS U1774 ( .A(n3457), .A(n3457_n), .B(n2836), .B(n2836_n), .Y(n2837_n), .Y(n2837) );
 NAND2X1TS U1775 ( .A(n3025), .A(n3025_n), .B(n3227), .B(n3227_n), .Y(n2838_n), .Y(n2838) );
 NAND2X1TS U1776 ( .A(n2837), .A(n2837_n), .B(n2838), .B(n2838_n), .Y(n2839_n), .Y(n2839) );
 NOR2X1TS U1777 ( .A(n3320), .A(n3320_n), .B(n3011), .B(n3011_n), .Y(n2840_n), .Y(n2840) );
 NOR2X1TS U1778 ( .A(n2840), .A(n2840_n), .B(n2839), .B(n2839_n), .Y(n2841_n), .Y(n2841) );
 NAND2BX1TS U1779 ( .AN(n3412), .AN(n3412_n), .B(n2998), .B(n2998_n), .Y(n2842_n), .Y(n2842) );
 NAND2X1TS U1780 ( .A(n2841), .A(n2841_n), .B(n2842), .B(n2842_n), .Y(n2843_n), .Y(n2843) );
 NOR2X1TS U1781 ( .A(n2835), .A(n2835_n), .B(n2843), .B(n2843_n), .Y(n2844_n), .Y(n2844) );
 NOR2X1TS U1782 ( .A(n3723), .A(n3723_n), .B(n3724), .B(n3724_n), .Y(n2845_n), .Y(n2845) );
 NAND2X1TS U1783 ( .A(n2844), .A(n2844_n), .B(n2845), .B(n2845_n), .Y(n2846_n), .Y(n2846) );
 NOR2X1TS U1784 ( .A(n2832), .A(n2832_n), .B(n2846), .B(n2846_n), .Y(n2847_n), .Y(n2847) );
 NOR2X1TS U1785 ( .A(n3598), .A(n3598_n), .B(n3331), .B(n3331_n), .Y(n2848_n), .Y(n2848) );
 NAND2X1TS U1786 ( .A(n2847), .A(n2847_n), .B(n2848), .B(n2848_n), .Y(n2849_n), .Y(n2849) );
 NOR2BX1TS U1787 ( .AN(n3620), .AN(n3620_n), .B(n2849), .B(n2849_n), .Y(n2850_n), .Y(n2850) );
 NAND2X1TS U1788 ( .A(n3124), .A(n3124_n), .B(n2850), .B(n2850_n), .Y(d[0]_n), .Y(d[0]) );
 NOR2BX1TS U1789 ( .AN(n3377), .AN(n3377_n), .B(n3164), .B(n3164_n), .Y(n2851_n), .Y(n2851) );
 NOR2X1TS U1790 ( .A(n3309), .A(n3309_n), .B(n3386), .B(n3386_n), .Y(n2852_n), .Y(n2852) );
 NAND2X1TS U1791 ( .A(n2851), .A(n2851_n), .B(n2852), .B(n2852_n), .Y(n2853_n), .Y(n2853) );
 NAND2X1TS U1792 ( .A(n3061), .A(n3061_n), .B(n3393), .B(n3393_n), .Y(n2854_n), .Y(n2854) );
 NAND2X1TS U1793 ( .A(n3588), .A(n3588_n), .B(n2854), .B(n2854_n), .Y(n2855_n), .Y(n2855) );
 NOR2X1TS U1794 ( .A(n2853), .A(n2853_n), .B(n2855), .B(n2855_n), .Y(n2856_n), .Y(n2856) );
 NOR2X1TS U1795 ( .A(n3281), .A(n3281_n), .B(n3587), .B(n3587_n), .Y(n2857_n), .Y(n2857) );
 NAND2X1TS U1796 ( .A(n2856), .A(n2856_n), .B(n2857), .B(n2857_n), .Y(n2858_n), .Y(n2858) );
 NAND2X1TS U1797 ( .A(n3414), .A(n3414_n), .B(n3416), .B(n3416_n), .Y(n2859_n), .Y(n2859) );
 NAND2X1TS U1798 ( .A(n3415), .A(n3415_n), .B(n3413), .B(n3413_n), .Y(n2860_n), .Y(n2860) );
 NOR2X1TS U1799 ( .A(n3016), .A(n3016_n), .B(n3412), .B(n3412_n), .Y(n2861_n), .Y(n2861) );
 NOR2X1TS U1800 ( .A(n3054), .A(n3054_n), .B(n3337), .B(n3337_n), .Y(n2862_n), .Y(n2862) );
 NOR2X1TS U1801 ( .A(n2859), .A(n2859_n), .B(n2860), .B(n2860_n), .Y(n2863_n), .Y(n2863) );
 NOR2X1TS U1802 ( .A(n2861), .A(n2861_n), .B(n2862), .B(n2862_n), .Y(n2864_n), .Y(n2864) );
 NAND2X1TS U1803 ( .A(n2863), .A(n2863_n), .B(n2864), .B(n2864_n), .Y(n2865_n), .Y(n2865) );
 NOR2X1TS U1804 ( .A(n3027), .A(n3027_n), .B(n3064), .B(n3064_n), .Y(n2866_n), .Y(n2866) );
 NOR2X1TS U1805 ( .A(n2954), .A(n2954_n), .B(n2866), .B(n2866_n), .Y(n2867_n), .Y(n2867) );
 NOR2X1TS U1806 ( .A(n2858), .A(n2858_n), .B(n2865), .B(n2865_n), .Y(n2868_n), .Y(n2868) );
 NOR2X1TS U1807 ( .A(n3411), .A(n3411_n), .B(n2867), .B(n2867_n), .Y(n2869_n), .Y(n2869) );
 NAND2X1TS U1808 ( .A(n2868), .A(n2868_n), .B(n2869), .B(n2869_n), .Y(d[2]_n), .Y(d[2]) );
 NAND2X1TS U1809 ( .A(n3064), .A(n3064_n), .B(n2969), .B(n2969_n), .Y(n2870_n), .Y(n2870) );
 NAND2X1TS U1810 ( .A(n3313), .A(n3313_n), .B(n2870), .B(n2870_n), .Y(n2871_n), .Y(n2871) );
 NAND2X1TS U1811 ( .A(n3216), .A(n3216_n), .B(n3314), .B(n3314_n), .Y(n2872_n), .Y(n2872) );
 NAND2X1TS U1812 ( .A(n2942), .A(n2942_n), .B(n3315), .B(n3315_n), .Y(n2873_n), .Y(n2873) );
 NAND2X1TS U1813 ( .A(n2872), .A(n2872_n), .B(n2873), .B(n2873_n), .Y(n2874_n), .Y(n2874) );
 NAND2X1TS U1814 ( .A(n3076), .A(n3076_n), .B(n3318), .B(n3318_n), .Y(n2875_n), .Y(n2875) );
 NAND2X1TS U1815 ( .A(n3317), .A(n3317_n), .B(n2875), .B(n2875_n), .Y(n2876_n), .Y(n2876) );
 NAND2X1TS U1816 ( .A(n3322), .A(n3322_n), .B(n3078), .B(n3078_n), .Y(n2877_n), .Y(n2877) );
 NAND2X1TS U1817 ( .A(n3018), .A(n3018_n), .B(n3250), .B(n3250_n), .Y(n2878_n), .Y(n2878) );
 NAND2X1TS U1818 ( .A(n2877), .A(n2877_n), .B(n2878), .B(n2878_n), .Y(n2879_n), .Y(n2879) );
 NOR2X1TS U1819 ( .A(n2871), .A(n2871_n), .B(n2874), .B(n2874_n), .Y(n2880_n), .Y(n2880) );
 NOR2X1TS U1820 ( .A(n2876), .A(n2876_n), .B(n2879), .B(n2879_n), .Y(n2881_n), .Y(n2881) );
 NAND2X1TS U1821 ( .A(n2880), .A(n2880_n), .B(n2881), .B(n2881_n), .Y(n2882_n), .Y(n2882) );
 OR2X1TS U1822 ( .A(n3385), .A(n3385_n), .B(n3386), .B(n3386_n), .Y(n2883_n), .Y(n2883) );
 NAND2X1TS U1823 ( .A(n3384), .A(n3384_n), .B(n3383), .B(n3383_n), .Y(n2884_n), .Y(n2884) );
 NOR2X1TS U1824 ( .A(n2883), .A(n2883_n), .B(n2884), .B(n2884_n), .Y(n2885_n), .Y(n2885) );
 NOR2X1TS U1825 ( .A(n3281), .A(n3281_n), .B(n3270), .B(n3270_n), .Y(n2886_n), .Y(n2886) );
 NAND2X1TS U1826 ( .A(n2885), .A(n2885_n), .B(n2886), .B(n2886_n), .Y(n2887_n), .Y(n2887) );
 NOR2X1TS U1827 ( .A(n2882), .A(n2882_n), .B(n2887), .B(n2887_n), .Y(n2888_n), .Y(n2888) );
 NAND2X1TS U1828 ( .A(n3191), .A(n3191_n), .B(n2888), .B(n2888_n), .Y(d[3]_n), .Y(d[3]) );
 NAND2BX1TS U1829 ( .AN(n3185), .AN(n3185_n), .B(n3184), .B(n3184_n), .Y(n3150_n), .Y(n3150) );
 NOR2X1TS U1830 ( .A(n3218), .A(n3218_n), .B(n3264), .B(n3264_n), .Y(n2889_n), .Y(n2889) );
 NAND2BX1TS U1831 ( .AN(n3311), .AN(n3311_n), .B(n3312), .B(n3312_n), .Y(n2890_n), .Y(n2890) );
 NOR2X1TS U1832 ( .A(n2889), .A(n2889_n), .B(n2890), .B(n2890_n), .Y(n2891_n), .Y(n2891) );
 NAND2X1TS U1833 ( .A(n3310), .A(n3310_n), .B(n2891), .B(n2891_n), .Y(n2892_n), .Y(n2892) );
 NOR2X1TS U1834 ( .A(n3274), .A(n3274_n), .B(n3275), .B(n3275_n), .Y(n2893_n), .Y(n2893) );
 NOR2X1TS U1835 ( .A(n3278), .A(n3278_n), .B(n3279), .B(n3279_n), .Y(n2894_n), .Y(n2894) );
 NAND2X1TS U1836 ( .A(n2893), .A(n2893_n), .B(n2894), .B(n2894_n), .Y(n2895_n), .Y(n2895) );
 NAND2X1TS U1837 ( .A(n3077), .A(n3077_n), .B(n3271), .B(n3271_n), .Y(n2896_n), .Y(n2896) );
 NAND2X1TS U1838 ( .A(n2973), .A(n2973_n), .B(n3008), .B(n3008_n), .Y(n2897_n), .Y(n2897) );
 NAND2X1TS U1839 ( .A(n2896), .A(n2896_n), .B(n2897), .B(n2897_n), .Y(n2898_n), .Y(n2898) );
 NOR2X1TS U1840 ( .A(n3149), .A(n3149_n), .B(n2935), .B(n2935_n), .Y(n2899_n), .Y(n2899) );
 AND2X1TS U1841 ( .A(n2968), .A(n2968_n), .B(n3272), .B(n3272_n), .Y(n2900_n), .Y(n2900) );
 NOR2X1TS U1842 ( .A(n2895), .A(n2895_n), .B(n2898), .B(n2898_n), .Y(n2901_n), .Y(n2901) );
 NOR2X1TS U1843 ( .A(n2899), .A(n2899_n), .B(n2900), .B(n2900_n), .Y(n2902_n), .Y(n2902) );
 NAND2X1TS U1844 ( .A(n2901), .A(n2901_n), .B(n2902), .B(n2902_n), .Y(n2903_n), .Y(n2903) );
 NOR2X1TS U1845 ( .A(n2892), .A(n2892_n), .B(n2903), .B(n2903_n), .Y(n2904_n), .Y(n2904) );
 NOR2X1TS U1846 ( .A(n3270), .A(n3270_n), .B(n3273), .B(n3273_n), .Y(n2905_n), .Y(n2905) );
 NAND2X1TS U1847 ( .A(n2904), .A(n2904_n), .B(n2905), .B(n2905_n), .Y(n2906_n), .Y(n2906) );
 NOR2X1TS U1848 ( .A(n3309), .A(n3309_n), .B(n2906), .B(n2906_n), .Y(n2907_n), .Y(n2907) );
 NAND2X1TS U1849 ( .A(n3162), .A(n3162_n), .B(n2907), .B(n2907_n), .Y(d[4]_n), .Y(d[4]) );
 OR2X2TS U1850 ( .A(n3804), .A(n3804_n), .B(n3858), .B(n3858_n), .Y(n2908_n), .Y(n2908) );
 OR2X2TS U1851 ( .A(n2999), .A(n2999_n), .B(n3802), .B(n3802_n), .Y(n2909_n), .Y(n2909) );
 OR2X2TS U1852 ( .A(n3120), .A(n3120_n), .B(n3510), .B(n3510_n), .Y(n2910_n), .Y(n2910) );
 AND2X2TS U1853 ( .A(n3104), .A(n3104_n), .B(n3871), .B(n3871_n), .Y(n2911_n), .Y(n2911) );
 NAND2X1TS U1854 ( .A(n3108), .A(n3108_n), .B(n3877), .B(n3877_n), .Y(n2912_n), .Y(n2912) );
 AND2X2TS U1855 ( .A(n2984), .A(n2984_n), .B(n2979), .B(n2979_n), .Y(n2913_n), .Y(n2913) );
 AND2X2TS U1856 ( .A(n3828), .A(n3828_n), .B(n3863), .B(n3863_n), .Y(n2914_n), .Y(n2914) );
 AND2X2TS U1857 ( .A(n2911), .A(n2911_n), .B(n3094), .B(n3094_n), .Y(n2915_n), .Y(n2915) );
 OR2X2TS U1858 ( .A(n3804), .A(n3804_n), .B(n2962), .B(n2962_n), .Y(n2916_n), .Y(n2916) );
 OR2X2TS U1859 ( .A(n3078), .A(n3078_n), .B(n3007), .B(n3007_n), .Y(n2917_n), .Y(n2917) );
 OR2X2TS U1860 ( .A(n3111), .A(n3111_n), .B(n3228), .B(n3228_n), .Y(n2918_n), .Y(n2918) );
 AND2X2TS U1861 ( .A(n3721), .A(n3721_n), .B(n3093), .B(n3093_n), .Y(n2919_n), .Y(n2919) );
 AND2X2TS U1862 ( .A(n2996), .A(n2996_n), .B(n3096), .B(n3096_n), .Y(n2920_n), .Y(n2920) );
 OR2X2TS U1863 ( .A(n3122), .A(n3122_n), .B(n3087), .B(n3087_n), .Y(n2921_n), .Y(n2921) );
 AND2X2TS U1864 ( .A(n3000), .A(n3000_n), .B(n3863), .B(n3863_n), .Y(n2922_n), .Y(n2922) );
 OR2X2TS U1865 ( .A(n3095), .A(n3095_n), .B(n3037), .B(n3037_n), .Y(n2923_n), .Y(n2923) );
 AND2X2TS U1866 ( .A(n2944), .A(n2944_n), .B(n3096), .B(n3096_n), .Y(n2924_n), .Y(n2924) );
 OR2X2TS U1867 ( .A(n3093), .A(n3093_n), .B(n3090), .B(n3090_n), .Y(n2925_n), .Y(n2925) );
 AND2X2TS U1868 ( .A(n2974), .A(n2974_n), .B(n3030), .B(n3030_n), .Y(n2926_n), .Y(n2926) );
 OR2X2TS U1869 ( .A(n3117), .A(n3117_n), .B(n3858), .B(n3858_n), .Y(n2927_n), .Y(n2927) );
 OR2X2TS U1870 ( .A(n3118), .A(n3118_n), .B(n3435), .B(n3435_n), .Y(n2928_n), .Y(n2928) );
 OR2X2TS U1871 ( .A(n3117), .A(n3117_n), .B(n3812), .B(n3812_n), .Y(n2929_n), .Y(n2929) );
 OR2X2TS U1872 ( .A(n3030), .A(n3030_n), .B(n3713), .B(n3713_n), .Y(n2930_n), .Y(n2930) );
 AND2X2TS U1873 ( .A(n3078), .A(n3078_n), .B(n3093), .B(n3093_n), .Y(n2931_n), .Y(n2931) );
 AND2X2TS U1874 ( .A(n2978), .A(n2978_n), .B(n3007), .B(n3007_n), .Y(n2932_n), .Y(n2932) );
 INVXLTS U1875 ( .A(n2916), .A(n2916_n), .Y(n2933_n), .Y(n2933) );
 INVXLTS U1876 ( .A(n2916), .A(n2916_n), .Y(n2934_n), .Y(n2934) );
 INVXLTS U1877 ( .A(n2917), .A(n2917_n), .Y(n2935_n), .Y(n2935) );
 INVXLTS U1878 ( .A(n2917), .A(n2917_n), .Y(n2936_n), .Y(n2936) );
 INVXLTS U1879 ( .A(n3298), .A(n3298_n), .Y(n2937_n), .Y(n2937) );
 INVXLTS U1880 ( .A(n3298), .A(n3298_n), .Y(n2938_n), .Y(n2938) );
 INVXLTS U1881 ( .A(n3417), .A(n3417_n), .Y(n2939_n), .Y(n2939) );
 INVXLTS U1882 ( .A(n3417), .A(n3417_n), .Y(n2940_n), .Y(n2940) );
 INVXLTS U1883 ( .A(n3257), .A(n3257_n), .Y(n2941_n), .Y(n2941) );
 INVXLTS U1884 ( .A(n2941), .A(n2941_n), .Y(n2942_n), .Y(n2942) );
 INVXLTS U1885 ( .A(n3393), .A(n3393_n), .Y(n2943_n), .Y(n2943) );
 INVXLTS U1886 ( .A(n2943), .A(n2943_n), .Y(n2944_n), .Y(n2944) );
 INVXLTS U1887 ( .A(n2920), .A(n2920_n), .Y(n2945_n), .Y(n2945) );
 INVXLTS U1888 ( .A(n2920), .A(n2920_n), .Y(n2946_n), .Y(n2946) );
 INVXLTS U1889 ( .A(n3319), .A(n3319_n), .Y(n2947_n), .Y(n2947) );
 INVXLTS U1890 ( .A(n3319), .A(n3319_n), .Y(n2948_n), .Y(n2948) );
 INVXLTS U1891 ( .A(n3215), .A(n3215_n), .Y(n2949_n), .Y(n2949) );
 INVXLTS U1892 ( .A(n2949), .A(n2949_n), .Y(n2950_n), .Y(n2950) );
 INVXLTS U1893 ( .A(n3457), .A(n3457_n), .Y(n2951_n), .Y(n2951) );
 INVXLTS U1894 ( .A(n2951), .A(n2951_n), .Y(n2952_n), .Y(n2952) );
 INVXLTS U1895 ( .A(n2913), .A(n2913_n), .Y(n2953_n), .Y(n2953) );
 INVXLTS U1896 ( .A(n2913), .A(n2913_n), .Y(n2954_n), .Y(n2954) );
 INVXLTS U1897 ( .A(n3465), .A(n3465_n), .Y(n2955_n), .Y(n2955) );
 INVXLTS U1898 ( .A(n2955), .A(n2955_n), .Y(n2956_n), .Y(n2956) );
 INVXLTS U1899 ( .A(n2930), .A(n2930_n), .Y(n2957_n), .Y(n2957) );
 INVXLTS U1900 ( .A(n2930), .A(n2930_n), .Y(n2958_n), .Y(n2958) );
 INVXLTS U1901 ( .A(n3119), .A(n3119_n), .Y(n2959_n), .Y(n2959) );
 INVXLTS U1902 ( .A(n2931), .A(n2931_n), .Y(n2960_n), .Y(n2960) );
 INVXLTS U1903 ( .A(n2931), .A(n2931_n), .Y(n2961_n), .Y(n2961) );
 INVXLTS U1904 ( .A(n2919), .A(n2919_n), .Y(n2962_n), .Y(n2962) );
 INVXLTS U1905 ( .A(n2919), .A(n2919_n), .Y(n2963_n), .Y(n2963) );
 INVXLTS U1906 ( .A(n2928), .A(n2928_n), .Y(n2964_n), .Y(n2964) );
 INVXLTS U1907 ( .A(n2928), .A(n2928_n), .Y(n2965_n), .Y(n2965) );
 INVXLTS U1908 ( .A(n2929), .A(n2929_n), .Y(n2966_n), .Y(n2966) );
 INVXLTS U1909 ( .A(n2929), .A(n2929_n), .Y(n2967_n), .Y(n2967) );
 INVXLTS U1910 ( .A(n3768), .A(n3768_n), .Y(n2968_n), .Y(n2968) );
 INVXLTS U1911 ( .A(n3768), .A(n3768_n), .Y(n2969_n), .Y(n2969) );
 INVXLTS U1912 ( .A(n3721), .A(n3721_n), .Y(n2970_n), .Y(n2970) );
 INVXLTS U1913 ( .A(n2970), .A(n2970_n), .Y(n2971_n), .Y(n2971) );
 INVXLTS U1914 ( .A(n3140), .A(n3140_n), .Y(n2972_n), .Y(n2972) );
 INVXLTS U1915 ( .A(n2972), .A(n2972_n), .Y(n2973_n), .Y(n2973) );
 INVXLTS U1916 ( .A(n2927), .A(n2927_n), .Y(n2974_n), .Y(n2974) );
 INVXLTS U1917 ( .A(n2927), .A(n2927_n), .Y(n2975_n), .Y(n2975) );
 INVXLTS U1918 ( .A(n3121), .A(n3121_n), .Y(n2976_n), .Y(n2976) );
 INVXLTS U1919 ( .A(n2976), .A(n2976_n), .Y(n2977_n), .Y(n2977) );
 INVXLTS U1920 ( .A(n3093), .A(n3093_n), .Y(n2978_n), .Y(n2978) );
 INVXLTS U1921 ( .A(n2978), .A(n2978_n), .Y(n2979_n), .Y(n2979) );
 INVXLTS U1922 ( .A(n3276), .A(n3276_n), .Y(n2980_n), .Y(n2980) );
 INVXLTS U1923 ( .A(n2980), .A(n2980_n), .Y(n2981_n), .Y(n2981) );
 INVXLTS U1924 ( .A(n3322), .A(n3322_n), .Y(n2982_n), .Y(n2982) );
 INVXLTS U1925 ( .A(n2982), .A(n2982_n), .Y(n2983_n), .Y(n2983) );
 INVXLTS U1926 ( .A(n3235), .A(n3235_n), .Y(n2984_n), .Y(n2984) );
 INVXLTS U1927 ( .A(n3235), .A(n3235_n), .Y(n2985_n), .Y(n2985) );
 INVXLTS U1928 ( .A(n3307), .A(n3307_n), .Y(n2986_n), .Y(n2986) );
 INVXLTS U1929 ( .A(n3307), .A(n3307_n), .Y(n2987_n), .Y(n2987) );
 INVXLTS U1930 ( .A(n2923), .A(n2923_n), .Y(n2988_n), .Y(n2988) );
 INVXLTS U1931 ( .A(n2923), .A(n2923_n), .Y(n2989_n), .Y(n2989) );
 INVXLTS U1932 ( .A(n2921), .A(n2921_n), .Y(n2990_n), .Y(n2990) );
 INVXLTS U1933 ( .A(n2921), .A(n2921_n), .Y(n2991_n), .Y(n2991) );
 INVXLTS U1934 ( .A(n3216), .A(n3216_n), .Y(n2992_n), .Y(n2992) );
 INVXLTS U1935 ( .A(n2992), .A(n2992_n), .Y(n2993_n), .Y(n2993) );
 INVXLTS U1936 ( .A(n2912), .A(n2912_n), .Y(n2994_n), .Y(n2994) );
 INVXLTS U1937 ( .A(n2912), .A(n2912_n), .Y(n2995_n), .Y(n2995) );
 INVXLTS U1938 ( .A(n3764), .A(n3764_n), .Y(n2996_n), .Y(n2996) );
 INVXLTS U1939 ( .A(n2925), .A(n2925_n), .Y(n2997_n), .Y(n2997) );
 INVXLTS U1940 ( .A(n2925), .A(n2925_n), .Y(n2998_n), .Y(n2998) );
 INVXLTS U1941 ( .A(n3184), .A(n3184_n), .Y(n2999_n), .Y(n2999) );
 INVXLTS U1942 ( .A(n2999), .A(n2999_n), .Y(n3000_n), .Y(n3000) );
 INVXLTS U1943 ( .A(n3597), .A(n3597_n), .Y(n3001_n), .Y(n3001) );
 INVXLTS U1944 ( .A(n3001), .A(n3001_n), .Y(n3002_n), .Y(n3002) );
 INVXLTS U1945 ( .A(n3174), .A(n3174_n), .Y(n3003_n), .Y(n3003) );
 INVXLTS U1946 ( .A(n3003), .A(n3003_n), .Y(n3004_n), .Y(n3004) );
 INVXLTS U1947 ( .A(n2926), .A(n2926_n), .Y(n3005_n), .Y(n3005) );
 INVXLTS U1948 ( .A(n2926), .A(n2926_n), .Y(n3006_n), .Y(n3006) );
 INVXLTS U1949 ( .A(n3316), .A(n3316_n), .Y(n3007_n), .Y(n3007) );
 INVXLTS U1950 ( .A(n3316), .A(n3316_n), .Y(n3008_n), .Y(n3008) );
 INVXLTS U1951 ( .A(n2924), .A(n2924_n), .Y(n3009_n), .Y(n3009) );
 INVXLTS U1952 ( .A(n2924), .A(n2924_n), .Y(n3010_n), .Y(n3010) );
 INVXLTS U1953 ( .A(n3233), .A(n3233_n), .Y(n3011_n), .Y(n3011) );
 INVXLTS U1954 ( .A(n3233), .A(n3233_n), .Y(n3012_n), .Y(n3012) );
 INVXLTS U1955 ( .A(n2915), .A(n2915_n), .Y(n3013_n), .Y(n3013) );
 INVXLTS U1956 ( .A(n2915), .A(n2915_n), .Y(n3014_n), .Y(n3014) );
 INVXLTS U1957 ( .A(n2932), .A(n2932_n), .Y(n3015_n), .Y(n3015) );
 INVXLTS U1958 ( .A(n2932), .A(n2932_n), .Y(n3016_n), .Y(n3016) );
 INVXLTS U1959 ( .A(n2986), .A(n2986_n), .Y(n3017_n), .Y(n3017) );
 INVXLTS U1960 ( .A(n2987), .A(n2987_n), .Y(n3018_n), .Y(n3018) );
 INVXLTS U1961 ( .A(n2922), .A(n2922_n), .Y(n3019_n), .Y(n3019) );
 INVXLTS U1962 ( .A(n2922), .A(n2922_n), .Y(n3020_n), .Y(n3020) );
 INVXLTS U1963 ( .A(n2918), .A(n2918_n), .Y(n3021_n), .Y(n3021) );
 INVXLTS U1964 ( .A(n2918), .A(n2918_n), .Y(n3022_n), .Y(n3022) );
 INVXLTS U1965 ( .A(n2914), .A(n2914_n), .Y(n3023_n), .Y(n3023) );
 INVXLTS U1966 ( .A(n2914), .A(n2914_n), .Y(n3024_n), .Y(n3024) );
 INVXLTS U1967 ( .A(n3175), .A(n3175_n), .Y(n3025_n), .Y(n3025) );
 INVXLTS U1968 ( .A(n3175), .A(n3175_n), .Y(n3026_n), .Y(n3026) );
 INVXLTS U1969 ( .A(n3173), .A(n3173_n), .Y(n3027_n), .Y(n3027) );
 INVXLTS U1970 ( .A(n3173), .A(n3173_n), .Y(n3028_n), .Y(n3028) );
 INVXLTS U1971 ( .A(n3113), .A(n3113_n), .Y(n3029_n), .Y(n3029) );
 INVXLTS U1972 ( .A(n3114), .A(n3114_n), .Y(n3030_n), .Y(n3030) );
 INVXLTS U1973 ( .A(n3308), .A(n3308_n), .Y(n3031_n), .Y(n3031) );
 INVXLTS U1974 ( .A(n3031), .A(n3031_n), .Y(n3032_n), .Y(n3032) );
 INVXLTS U1975 ( .A(n3345), .A(n3345_n), .Y(n3033_n), .Y(n3033) );
 INVXLTS U1976 ( .A(n3033), .A(n3033_n), .Y(n3034_n), .Y(n3034) );
 INVXLTS U1977 ( .A(n3033), .A(n3033_n), .Y(n3035_n), .Y(n3035) );
 INVXLTS U1978 ( .A(n3265), .A(n3265_n), .Y(n3036_n), .Y(n3036) );
 INVXLTS U1979 ( .A(n3036), .A(n3036_n), .Y(n3037_n), .Y(n3037) );
 INVXLTS U1980 ( .A(n3036), .A(n3036_n), .Y(n3038_n), .Y(n3038) );
 INVXLTS U1981 ( .A(n2939), .A(n2939_n), .Y(n3039_n), .Y(n3039) );
 INVXLTS U1982 ( .A(n2940), .A(n2940_n), .Y(n3040_n), .Y(n3040) );
 INVXLTS U1983 ( .A(n2910), .A(n2910_n), .Y(n3041_n), .Y(n3041) );
 INVXLTS U1984 ( .A(n2910), .A(n2910_n), .Y(n3043_n), .Y(n3043) );
 INVXLTS U1985 ( .A(n2910), .A(n2910_n), .Y(n3042_n), .Y(n3042) );
 INVXLTS U1986 ( .A(n2937), .A(n2937_n), .Y(n3044_n), .Y(n3044) );
 INVXLTS U1987 ( .A(n2938), .A(n2938_n), .Y(n3045_n), .Y(n3045) );
 INVXLTS U1988 ( .A(n3173), .A(n3173_n), .Y(n3046_n), .Y(n3046) );
 INVXLTS U1989 ( .A(n3046), .A(n3046_n), .Y(n3047_n), .Y(n3047) );
 INVXLTS U1990 ( .A(n3046), .A(n3046_n), .Y(n3048_n), .Y(n3048) );
 INVXLTS U1991 ( .A(n2947), .A(n2947_n), .Y(n3049_n), .Y(n3049) );
 INVXLTS U1992 ( .A(n2948), .A(n2948_n), .Y(n3050_n), .Y(n3050) );
 INVXLTS U1993 ( .A(n2994), .A(n2994_n), .Y(n3051_n), .Y(n3051) );
 INVXLTS U1994 ( .A(n2995), .A(n2995_n), .Y(n3052_n), .Y(n3052) );
 INVXLTS U1995 ( .A(n2911), .A(n2911_n), .Y(n3053_n), .Y(n3053) );
 INVXLTS U1996 ( .A(n2911), .A(n2911_n), .Y(n3055_n), .Y(n3055) );
 INVXLTS U1997 ( .A(n2911), .A(n2911_n), .Y(n3054_n), .Y(n3054) );
 INVXLTS U1998 ( .A(n3175), .A(n3175_n), .Y(n3056_n), .Y(n3056) );
 INVXLTS U1999 ( .A(n3056), .A(n3056_n), .Y(n3057_n), .Y(n3057) );
 INVXLTS U2000 ( .A(n3056), .A(n3056_n), .Y(n3059_n), .Y(n3059) );
 INVXLTS U2001 ( .A(n3056), .A(n3056_n), .Y(n3058_n), .Y(n3058) );
 INVXLTS U2002 ( .A(n2908), .A(n2908_n), .Y(n3060_n), .Y(n3060) );
 INVXLTS U2003 ( .A(n2908), .A(n2908_n), .Y(n3062_n), .Y(n3062) );
 INVXLTS U2004 ( .A(n2908), .A(n2908_n), .Y(n3061_n), .Y(n3061) );
 INVXLTS U2005 ( .A(n3146), .A(n3146_n), .Y(n3063_n), .Y(n3063) );
 INVXLTS U2006 ( .A(n3063), .A(n3063_n), .Y(n3064_n), .Y(n3064) );
 INVXLTS U2007 ( .A(n3063), .A(n3063_n), .Y(n3065_n), .Y(n3065) );
 INVXLTS U2008 ( .A(n2909), .A(n2909_n), .Y(n3066_n), .Y(n3066) );
 INVXLTS U2009 ( .A(n2909), .A(n2909_n), .Y(n3068_n), .Y(n3068) );
 INVXLTS U2010 ( .A(n2909), .A(n2909_n), .Y(n3067_n), .Y(n3067) );
 INVXLTS U2011 ( .A(n2924), .A(n2924_n), .Y(n3069_n), .Y(n3069) );
 INVXLTS U2012 ( .A(n3069), .A(n3069_n), .Y(n3070_n), .Y(n3070) );
 INVXLTS U2013 ( .A(n3069), .A(n3069_n), .Y(n3072_n), .Y(n3072) );
 INVXLTS U2014 ( .A(n3069), .A(n3069_n), .Y(n3071_n), .Y(n3071) );
 INVXLTS U2015 ( .A(n3233), .A(n3233_n), .Y(n3073_n), .Y(n3073) );
 INVXLTS U2016 ( .A(n3073), .A(n3073_n), .Y(n3074_n), .Y(n3074) );
 INVXLTS U2017 ( .A(n3073), .A(n3073_n), .Y(n3076_n), .Y(n3076) );
 INVXLTS U2018 ( .A(n3073), .A(n3073_n), .Y(n3075_n), .Y(n3075) );
 INVXLTS U2019 ( .A(n3265), .A(n3265_n), .Y(n3077_n), .Y(n3077) );
 INVXLTS U2020 ( .A(n3265), .A(n3265_n), .Y(n3079_n), .Y(n3079) );
 INVXLTS U2021 ( .A(n3265), .A(n3265_n), .Y(n3078_n), .Y(n3078) );
 INVXLTS U2022 ( .A(n2922), .A(n2922_n), .Y(n3080_n), .Y(n3080) );
 INVXLTS U2023 ( .A(n3080), .A(n3080_n), .Y(n3081_n), .Y(n3081) );
 INVXLTS U2024 ( .A(n3080), .A(n3080_n), .Y(n3083_n), .Y(n3083) );
 INVXLTS U2025 ( .A(n3080), .A(n3080_n), .Y(n3082_n), .Y(n3082) );
 INVXLTS U2026 ( .A(n3316), .A(n3316_n), .Y(n3084_n), .Y(n3084) );
 INVXLTS U2027 ( .A(n3084), .A(n3084_n), .Y(n3085_n), .Y(n3085) );
 INVXLTS U2028 ( .A(n3084), .A(n3084_n), .Y(n3087_n), .Y(n3087) );
 INVXLTS U2029 ( .A(n3084), .A(n3084_n), .Y(n3086_n), .Y(n3086) );
 INVXLTS U2030 ( .A(n3155), .A(n3155_n), .Y(n3088_n), .Y(n3088) );
 INVXLTS U2031 ( .A(n3088), .A(n3088_n), .Y(n3089_n), .Y(n3089) );
 INVXLTS U2032 ( .A(n3088), .A(n3088_n), .Y(n3090_n), .Y(n3090) );
 INVXLTS U2033 ( .A(n3088), .A(n3088_n), .Y(n3091_n), .Y(n3091) );
 INVXLTS U2034 ( .A(n2976), .A(n2976_n), .Y(n3092_n), .Y(n3092) );
 INVXLTS U2035 ( .A(n3092), .A(n3092_n), .Y(n3093_n), .Y(n3093) );
 INVXLTS U2036 ( .A(n3092), .A(n3092_n), .Y(n3096_n), .Y(n3096) );
 INVXLTS U2037 ( .A(n3092), .A(n3092_n), .Y(n3094_n), .Y(n3094) );
 INVXLTS U2038 ( .A(n3092), .A(n3092_n), .Y(n3095_n), .Y(n3095) );
 INVXLTS U2039 ( .A(a[7]), .A(a[7]_n), .Y(n3097_n), .Y(n3097) );
 INVXLTS U2040 ( .A(n3097), .A(n3097_n), .Y(n3098_n), .Y(n3098) );
 INVXLTS U2041 ( .A(n3097), .A(n3097_n), .Y(n3099_n), .Y(n3099) );
 INVXLTS U2042 ( .A(a[6]), .A(a[6]_n), .Y(n3100_n), .Y(n3100) );
 INVXLTS U2043 ( .A(n3100), .A(n3100_n), .Y(n3101_n), .Y(n3101) );
 INVXLTS U2044 ( .A(n3100), .A(n3100_n), .Y(n3102_n), .Y(n3102) );
 INVXLTS U2045 ( .A(a[2]), .A(a[2]_n), .Y(n3103_n), .Y(n3103) );
 INVXLTS U2046 ( .A(n3103), .A(n3103_n), .Y(n3104_n), .Y(n3104) );
 INVXLTS U2047 ( .A(n3103), .A(n3103_n), .Y(n3105_n), .Y(n3105) );
 INVXLTS U2048 ( .A(a[3]), .A(a[3]_n), .Y(n3106_n), .Y(n3106) );
 INVXLTS U2049 ( .A(n3106), .A(n3106_n), .Y(n3107_n), .Y(n3107) );
 INVXLTS U2050 ( .A(n3106), .A(n3106_n), .Y(n3108_n), .Y(n3108) );
 INVXLTS U2051 ( .A(a[0]), .A(a[0]_n), .Y(n3109_n), .Y(n3109) );
 INVXLTS U2052 ( .A(n3109), .A(n3109_n), .Y(n3110_n), .Y(n3110) );
 INVXLTS U2053 ( .A(n3109), .A(n3109_n), .Y(n3111_n), .Y(n3111) );
 INVXLTS U2054 ( .A(a[5]), .A(a[5]_n), .Y(n3112_n), .Y(n3112) );
 INVXLTS U2055 ( .A(n3112), .A(n3112_n), .Y(n3113_n), .Y(n3113) );
 INVXLTS U2056 ( .A(n3112), .A(n3112_n), .Y(n3115_n), .Y(n3115) );
 INVXLTS U2057 ( .A(n3112), .A(n3112_n), .Y(n3114_n), .Y(n3114) );
 INVXLTS U2058 ( .A(a[4]), .A(a[4]_n), .Y(n3116_n), .Y(n3116) );
 INVXLTS U2059 ( .A(n3116), .A(n3116_n), .Y(n3117_n), .Y(n3117) );
 INVXLTS U2060 ( .A(n3116), .A(n3116_n), .Y(n3119_n), .Y(n3119) );
 INVXLTS U2061 ( .A(n3116), .A(n3116_n), .Y(n3118_n), .Y(n3118) );
 INVXLTS U2062 ( .A(a[1]), .A(a[1]_n), .Y(n3120_n), .Y(n3120) );
 INVXLTS U2063 ( .A(n3120), .A(n3120_n), .Y(n3121_n), .Y(n3121) );
 INVXLTS U2064 ( .A(n3120), .A(n3120_n), .Y(n3123_n), .Y(n3123) );
 INVXLTS U2065 ( .A(n3120), .A(n3120_n), .Y(n3122_n), .Y(n3122) );
 NOR2X1TS U2066 ( .A(n3025), .A(n3025_n), .B(n3018), .B(n3018_n), .Y(n3725_n), .Y(n3725) );
 NOR2X1TS U2067 ( .A(n3181), .A(n3181_n), .B(n3091), .B(n3091_n), .Y(n3176_n), .Y(n3176) );
 NOR2X1TS U2068 ( .A(n3182), .A(n3182_n), .B(n2957), .B(n2957_n), .Y(n3181_n), .Y(n3181) );
 NOR2X1TS U2069 ( .A(n3071), .A(n3071_n), .B(n3042), .B(n3042_n), .Y(n3252_n), .Y(n3252) );
 NOR2X1TS U2070 ( .A(n3090), .A(n3090_n), .B(n3291), .B(n3291_n), .Y(n3290_n), .Y(n3290) );
 NOR2X1TS U2071 ( .A(n3018), .A(n3018_n), .B(n3308), .B(n3308_n), .Y(n3305_n), .Y(n3305) );
 NOR2X1TS U2072 ( .A(n3089), .A(n3089_n), .B(n3156), .B(n3156_n), .Y(n3154_n), .Y(n3154) );
 NOR2X1TS U2073 ( .A(n3068), .A(n3068_n), .B(n3247), .B(n3247_n), .Y(n3825_n), .Y(n3825) );
 NOR2X1TS U2074 ( .A(n3083), .A(n3083_n), .B(n3247), .B(n3247_n), .Y(n3868_n), .Y(n3868) );
 NOR2X1TS U2075 ( .A(n3348), .A(n3348_n), .B(n3074), .B(n3074_n), .Y(n3346_n), .Y(n3346) );
 NOR2X1TS U2076 ( .A(n3022), .A(n3022_n), .B(n3079), .B(n3079_n), .Y(n3217_n), .Y(n3217) );
 NOR2X1TS U2077 ( .A(n2991), .A(n2991_n), .B(n3410), .B(n3410_n), .Y(n3409_n), .Y(n3409) );
 NOR2X1TS U2078 ( .A(n3091), .A(n3091_n), .B(n3443), .B(n3443_n), .Y(n3439_n), .Y(n3439) );
 NOR2X1TS U2079 ( .A(n2973), .A(n2973_n), .B(n2958), .B(n2958_n), .Y(n3463_n), .Y(n3463) );
 NOR2X1TS U2080 ( .A(n2993), .A(n2993_n), .B(n3044), .B(n3044_n), .Y(n3502_n), .Y(n3502) );
 NOR2X1TS U2081 ( .A(n3557), .A(n3557_n), .B(n3089), .B(n3089_n), .Y(n3552_n), .Y(n3552) );
 NOR2X1TS U2082 ( .A(n3322), .A(n3322_n), .B(n3257), .B(n3257_n), .Y(n3557_n), .Y(n3557) );
 NOR2X1TS U2083 ( .A(n3575), .A(n3575_n), .B(n3155), .B(n3155_n), .Y(n3574_n), .Y(n3574) );
 NOR2X1TS U2084 ( .A(n3081), .A(n3081_n), .B(n3068), .B(n3068_n), .Y(n3576_n), .Y(n3576) );
 NOR2X1TS U2085 ( .A(n3060), .A(n3060_n), .B(n3271), .B(n3271_n), .Y(n3606_n), .Y(n3606) );
 NOR2X1TS U2086 ( .A(n3041), .A(n3041_n), .B(n3375), .B(n3375_n), .Y(n3615_n), .Y(n3615) );
 NOR2X1TS U2087 ( .A(n2950), .A(n2950_n), .B(n3322), .B(n3322_n), .Y(n3756_n), .Y(n3756) );
 NOR2X1TS U2088 ( .A(n3179), .A(n3179_n), .B(n3045), .B(n3045_n), .Y(n3787_n), .Y(n3787) );
 NOR2X1TS U2089 ( .A(n3074), .A(n3074_n), .B(n2997), .B(n2997_n), .Y(n3634_n), .Y(n3634) );
 NOR2X1TS U2090 ( .A(n2983), .A(n2983_n), .B(n2933), .B(n2933_n), .Y(n3803_n), .Y(n3803) );
 NOR2X1TS U2091 ( .A(n3808), .A(n3808_n), .B(n3090), .B(n3090_n), .Y(n3807_n), .Y(n3807) );
 NOR2X1TS U2092 ( .A(n2974), .A(n2974_n), .B(n3215), .B(n3215_n), .Y(n3808_n), .Y(n3808) );
 INVX2TS U2093 ( .A(n3863), .A(n3863_n), .Y(n3804_n), .Y(n3804) );
 NOR2X1TS U2094 ( .A(n3066), .A(n3066_n), .B(n3044), .B(n3044_n), .Y(n3500_n), .Y(n3500) );
 NAND2X1TS U2095 ( .A(n3111), .A(n3111_n), .B(n3372), .B(n3372_n), .Y(n3316_n), .Y(n3316) );
 NOR2X1TS U2096 ( .A(n3725), .A(n3725_n), .B(n3013), .B(n3013_n), .Y(n3724_n), .Y(n3724) );
 NOR2X1TS U2097 ( .A(n3726), .A(n3726_n), .B(n3306), .B(n3306_n), .Y(n3723_n), .Y(n3723) );
 NOR2X1TS U2098 ( .A(n2965), .A(n2965_n), .B(n3198), .B(n3198_n), .Y(n3726_n), .Y(n3726) );
 OR2X2TS U2099 ( .A(n3159), .A(n3159_n), .B(n3160), .B(n3160_n), .Y(d[6]_n), .Y(d[6]) );
 NOR2X1TS U2100 ( .A(n3163), .A(n3163_n), .B(n3164), .B(n3164_n), .Y(n3161_n), .Y(n3161) );
 NOR2X1TS U2101 ( .A(n3167), .A(n3167_n), .B(n3168), .B(n3168_n), .Y(n3165_n), .Y(n3165) );
 NOR2X1TS U2102 ( .A(n3171), .A(n3171_n), .B(n3172), .B(n3172_n), .Y(n3170_n), .Y(n3170) );
 NOR2X1TS U2103 ( .A(n3173), .A(n3173_n), .B(n3174), .B(n3174_n), .Y(n3172_n), .Y(n3172) );
 NOR2X1TS U2104 ( .A(n3057), .A(n3057_n), .B(n2961), .B(n2961_n), .Y(n3171_n), .Y(n3171) );
 NOR2X1TS U2105 ( .A(n3176), .A(n3176_n), .B(n3177), .B(n3177_n), .Y(n3169_n), .Y(n3169) );
 NOR2X1TS U2106 ( .A(n3178), .A(n3178_n), .B(n3011), .B(n3011_n), .Y(n3177_n), .Y(n3177) );
 NOR2X1TS U2107 ( .A(n3179), .A(n3179_n), .B(n3180), .B(n3180_n), .Y(n3178_n), .Y(n3178) );
 NOR2X1TS U2108 ( .A(n3186), .A(n3186_n), .B(n3187), .B(n3187_n), .Y(n3183_n), .Y(n3183) );
 NOR2X1TS U2109 ( .A(n3192), .A(n3192_n), .B(n3193), .B(n3193_n), .Y(n3190_n), .Y(n3190) );
 NOR2X1TS U2110 ( .A(n3202), .A(n3202_n), .B(n3203), .B(n3203_n), .Y(n3201_n), .Y(n3201) );
 NOR2X1TS U2111 ( .A(n3238), .A(n3238_n), .B(n3239), .B(n3239_n), .Y(n3237_n), .Y(n3237) );
 NOR2X1TS U2112 ( .A(n3242), .A(n3242_n), .B(n3243), .B(n3243_n), .Y(n3240_n), .Y(n3240) );
 INVX2TS U2113 ( .A(n3252), .A(n3252_n), .Y(n3251_n), .Y(n3251) );
 NOR2X1TS U2114 ( .A(n3258), .A(n3258_n), .B(n3259), .B(n3259_n), .Y(n3253_n), .Y(n3253) );
 NOR2X1TS U2115 ( .A(n3266), .A(n3266_n), .B(n3267), .B(n3267_n), .Y(n3200_n), .Y(n3200) );
 NOR2X1TS U2116 ( .A(n3729), .A(n3729_n), .B(n3730), .B(n3730_n), .Y(n3269_n), .Y(n3269) );
 NOR2X1TS U2117 ( .A(n3732), .A(n3732_n), .B(n3733), .B(n3733_n), .Y(n3731_n), .Y(n3731) );
 NOR2X1TS U2118 ( .A(n3737), .A(n3737_n), .B(n3361), .B(n3361_n), .Y(n3194_n), .Y(n3194) );
 NOR2X1TS U2119 ( .A(n3738), .A(n3738_n), .B(n3086), .B(n3086_n), .Y(n3737_n), .Y(n3737) );
 AND2X2TS U2120 ( .A(n3741), .A(n3741_n), .B(n3742), .B(n3742_n), .Y(n3740_n), .Y(n3740) );
 NOR2X1TS U2121 ( .A(n3743), .A(n3743_n), .B(n3744), .B(n3744_n), .Y(n3741_n), .Y(n3741) );
 NOR2X1TS U2122 ( .A(n3252), .A(n3252_n), .B(n2987), .B(n2987_n), .Y(n3744_n), .Y(n3744) );
 NOR2X1TS U2123 ( .A(n3576), .A(n3576_n), .B(n3034), .B(n3034_n), .Y(n3743_n), .Y(n3743) );
 NOR2X1TS U2124 ( .A(n3745), .A(n3745_n), .B(n3746), .B(n3746_n), .Y(n3739_n), .Y(n3739) );
 NOR2X1TS U2125 ( .A(n3748), .A(n3748_n), .B(n3085), .B(n3085_n), .Y(n3745_n), .Y(n3745) );
 NOR2X1TS U2126 ( .A(n3419), .A(n3419_n), .B(n3449), .B(n3449_n), .Y(n3748_n), .Y(n3748) );
 NOR2X1TS U2127 ( .A(n2981), .A(n2981_n), .B(n3011), .B(n3011_n), .Y(n3275_n), .Y(n3275) );
 NOR2X1TS U2128 ( .A(n3277), .A(n3277_n), .B(n2937), .B(n2937_n), .Y(n3274_n), .Y(n3274) );
 NOR2X1TS U2129 ( .A(n3280), .A(n3280_n), .B(n2939), .B(n2939_n), .Y(n3279_n), .Y(n3279) );
 NOR2X1TS U2130 ( .A(n3054), .A(n3054_n), .B(n3174), .B(n3174_n), .Y(n3278_n), .Y(n3278) );
 NOR2X1TS U2131 ( .A(n3281), .A(n3281_n), .B(n3282), .B(n3282_n), .Y(n3162_n), .Y(n3162) );
 NOR2X1TS U2132 ( .A(n3285), .A(n3285_n), .B(n3286), .B(n3286_n), .Y(n3284_n), .Y(n3284) );
 NOR2X1TS U2133 ( .A(n3289), .A(n3289_n), .B(n3290), .B(n3290_n), .Y(n3287_n), .Y(n3287) );
 NOR2X1TS U2134 ( .A(n3292), .A(n3292_n), .B(n3012), .B(n3012_n), .Y(n3289_n), .Y(n3289) );
 NOR2X1TS U2135 ( .A(n3293), .A(n3293_n), .B(n3294), .B(n3294_n), .Y(n3283_n), .Y(n3283) );
 NOR2X1TS U2136 ( .A(n3303), .A(n3303_n), .B(n3304), .B(n3304_n), .Y(n3299_n), .Y(n3299) );
 NOR2X1TS U2137 ( .A(n2935), .A(n2935_n), .B(n3004), .B(n3004_n), .Y(n3304_n), .Y(n3304) );
 NOR2X1TS U2138 ( .A(n3305), .A(n3305_n), .B(n3306), .B(n3306_n), .Y(n3303_n), .Y(n3303) );
 NOR2X1TS U2139 ( .A(n3126), .A(n3126_n), .B(n3127), .B(n3127_n), .Y(n3125_n), .Y(n3125) );
 NOR2X1TS U2140 ( .A(n3130), .A(n3130_n), .B(n3131), .B(n3131_n), .Y(n3129_n), .Y(n3129) );
 NOR2X1TS U2141 ( .A(n3134), .A(n3134_n), .B(n3135), .B(n3135_n), .Y(n3133_n), .Y(n3133) );
 NOR2X1TS U2142 ( .A(n3142), .A(n3142_n), .B(n3143), .B(n3143_n), .Y(n3132_n), .Y(n3132) );
 NOR2X1TS U2143 ( .A(n3153), .A(n3153_n), .B(n3154), .B(n3154_n), .Y(n3152_n), .Y(n3152) );
 NOR2X1TS U2144 ( .A(n3157), .A(n3157_n), .B(n3158), .B(n3158_n), .Y(n3151_n), .Y(n3151) );
 NOR2X1TS U2145 ( .A(n3024), .A(n3024_n), .B(n3015), .B(n3015_n), .Y(n3158_n), .Y(n3158) );
 NOR2X1TS U2146 ( .A(n3205), .A(n3205_n), .B(n3206), .B(n3206_n), .Y(n3128_n), .Y(n3128) );
 NOR2X1TS U2147 ( .A(n3209), .A(n3209_n), .B(n3210), .B(n3210_n), .Y(n3208_n), .Y(n3208) );
 NOR2X1TS U2148 ( .A(n3047), .A(n3047_n), .B(n2953), .B(n2953_n), .Y(n3209_n), .Y(n3209) );
 NOR2X1TS U2149 ( .A(n3211), .A(n3211_n), .B(n3212), .B(n3212_n), .Y(n3207_n), .Y(n3207) );
 NOR2X1TS U2150 ( .A(n3217), .A(n3217_n), .B(n3218), .B(n3218_n), .Y(n3211_n), .Y(n3211) );
 NOR2X1TS U2151 ( .A(n3221), .A(n3221_n), .B(n3222), .B(n3222_n), .Y(n3220_n), .Y(n3220) );
 NOR2X1TS U2152 ( .A(n3228), .A(n3228_n), .B(n2945), .B(n2945_n), .Y(n3221_n), .Y(n3221) );
 NOR2X1TS U2153 ( .A(n3229), .A(n3229_n), .B(n3230), .B(n3230_n), .Y(n3219_n), .Y(n3219) );
 NOR2X1TS U2154 ( .A(n3790), .A(n3790_n), .B(n3791), .B(n3791_n), .Y(n3124_n), .Y(n3124) );
 NOR2X1TS U2155 ( .A(n3815), .A(n3815_n), .B(n3816), .B(n3816_n), .Y(n3792_n), .Y(n3792) );
 NOR2X1TS U2156 ( .A(n3419), .A(n3419_n), .B(n3003), .B(n3003_n), .Y(n3256_n), .Y(n3256) );
 NOR2X1TS U2157 ( .A(n3820), .A(n3820_n), .B(n3821), .B(n3821_n), .Y(n3817_n), .Y(n3817) );
 NOR2X1TS U2158 ( .A(n3114), .A(n3114_n), .B(n3321), .B(n3321_n), .Y(n3823_n), .Y(n3823) );
 NOR2X1TS U2159 ( .A(n3825), .A(n3825_n), .B(n3277), .B(n3277_n), .Y(n3820_n), .Y(n3820) );
 NOR2X1TS U2160 ( .A(n3830), .A(n3830_n), .B(n3831), .B(n3831_n), .Y(n3826_n), .Y(n3826) );
 NOR2X1TS U2161 ( .A(n3638), .A(n3638_n), .B(n3664), .B(n3664_n), .Y(n3836_n), .Y(n3836) );
 NOR2X1TS U2162 ( .A(n3852), .A(n3852_n), .B(n3853), .B(n3853_n), .Y(n3236_n), .Y(n3236) );
 NOR2X1TS U2163 ( .A(n3856), .A(n3856_n), .B(n3857), .B(n3857_n), .Y(n3855_n), .Y(n3855) );
 NOR2X1TS U2164 ( .A(n2912), .A(n2912_n), .B(n3768), .B(n3768_n), .Y(n3857_n), .Y(n3857) );
 NOR2X1TS U2165 ( .A(n3038), .A(n3038_n), .B(n3291), .B(n3291_n), .Y(n3856_n), .Y(n3856) );
 NOR2X1TS U2166 ( .A(n3860), .A(n3860_n), .B(n3861), .B(n3861_n), .Y(n3854_n), .Y(n3854) );
 NOR2X1TS U2167 ( .A(n3435), .A(n3435_n), .B(n3829), .B(n3829_n), .Y(n3860_n), .Y(n3860) );
 NOR2X1TS U2168 ( .A(n3866), .A(n3866_n), .B(n3867), .B(n3867_n), .Y(n3865_n), .Y(n3865) );
 NOR2X1TS U2169 ( .A(n3868), .A(n3868_n), .B(n3010), .B(n3010_n), .Y(n3867_n), .Y(n3867) );
 NOR2X1TS U2170 ( .A(n3870), .A(n3870_n), .B(n3055), .B(n3055_n), .Y(n3866_n), .Y(n3866) );
 NOR2X1TS U2171 ( .A(n3402), .A(n3402_n), .B(n3872), .B(n3872_n), .Y(n3870_n), .Y(n3870) );
 NOR2X1TS U2172 ( .A(n3493), .A(n3493_n), .B(n3873), .B(n3873_n), .Y(n3864_n), .Y(n3864) );
 NOR2X1TS U2173 ( .A(n3112), .A(n3112_n), .B(n3321), .B(n3321_n), .Y(n3180_n), .Y(n3180) );
 INVX2TS U2174 ( .A(n3824), .A(n3824_n), .Y(n3321_n), .Y(n3321) );
 NOR2X1TS U2175 ( .A(n3323), .A(n3323_n), .B(n3324), .B(n3324_n), .Y(n3191_n), .Y(n3191) );
 NOR2X1TS U2176 ( .A(n3326), .A(n3326_n), .B(n3327), .B(n3327_n), .Y(n3310_n), .Y(n3310) );
 NOR2X1TS U2177 ( .A(n3330), .A(n3330_n), .B(n3331), .B(n3331_n), .Y(n3329_n), .Y(n3329) );
 NOR2X1TS U2178 ( .A(n3048), .A(n3048_n), .B(n3218), .B(n3218_n), .Y(n3331_n), .Y(n3331) );
 NOR2X1TS U2179 ( .A(n3332), .A(n3332_n), .B(n3333), .B(n3333_n), .Y(n3328_n), .Y(n3328) );
 NOR2X1TS U2180 ( .A(n3337), .A(n3337_n), .B(n3087), .B(n3087_n), .Y(n3332_n), .Y(n3332) );
 NOR2X1TS U2181 ( .A(n3340), .A(n3340_n), .B(n3341), .B(n3341_n), .Y(n3339_n), .Y(n3339) );
 NOR2X1TS U2182 ( .A(n3346), .A(n3346_n), .B(n3347), .B(n3347_n), .Y(n3340_n), .Y(n3340) );
 NOR2X1TS U2183 ( .A(n3353), .A(n3353_n), .B(n3354), .B(n3354_n), .Y(n3325_n), .Y(n3325) );
 INVX2TS U2184 ( .A(n3361), .A(n3361_n), .Y(n3358_n), .Y(n3358) );
 NOR2X1TS U2185 ( .A(n3364), .A(n3364_n), .B(n3365), .B(n3365_n), .Y(n3363_n), .Y(n3363) );
 NOR2X1TS U2186 ( .A(n3368), .A(n3368_n), .B(n3057), .B(n3057_n), .Y(n3364_n), .Y(n3364) );
 NOR2X1TS U2187 ( .A(n3369), .A(n3369_n), .B(n3370), .B(n3370_n), .Y(n3362_n), .Y(n3362) );
 NOR2X1TS U2188 ( .A(n3374), .A(n3374_n), .B(n2938), .B(n2938_n), .Y(n3369_n), .Y(n3369) );
 NOR2X1TS U2189 ( .A(n3375), .A(n3375_n), .B(n3376), .B(n3376_n), .Y(n3374_n), .Y(n3374) );
 NOR2X1TS U2190 ( .A(n3379), .A(n3379_n), .B(n3380), .B(n3380_n), .Y(n3378_n), .Y(n3378) );
 NOR2X1TS U2191 ( .A(n3006), .A(n3006_n), .B(n3038), .B(n3038_n), .Y(n3379_n), .Y(n3379) );
 NOR2X1TS U2192 ( .A(n3389), .A(n3389_n), .B(n3390), .B(n3390_n), .Y(n3388_n), .Y(n3388) );
 NOR2X1TS U2193 ( .A(n3210), .A(n3210_n), .B(n3397), .B(n3397_n), .Y(n3394_n), .Y(n3394) );
 NOR2X1TS U2194 ( .A(n3023), .A(n3023_n), .B(n3034), .B(n3034_n), .Y(n3397_n), .Y(n3397) );
 NOR2X1TS U2195 ( .A(n3090), .A(n3090_n), .B(n3149), .B(n3149_n), .Y(n3210_n), .Y(n3210) );
 NOR2X1TS U2196 ( .A(n3398), .A(n3398_n), .B(n3399), .B(n3399_n), .Y(n3387_n), .Y(n3387) );
 NOR2X1TS U2197 ( .A(n3407), .A(n3407_n), .B(n3408), .B(n3408_n), .Y(n3404_n), .Y(n3404) );
 NOR2X1TS U2198 ( .A(n3409), .A(n3409_n), .B(n2986), .B(n2986_n), .Y(n3408_n), .Y(n3408) );
 NOR2X1TS U2199 ( .A(n2936), .A(n2936_n), .B(n2979), .B(n2979_n), .Y(n3410_n), .Y(n3410) );
 NOR2X1TS U2200 ( .A(n3347), .A(n3347_n), .B(n3492), .B(n3492_n), .Y(n3411_n), .Y(n3411) );
 NOR2X1TS U2201 ( .A(n3392), .A(n3392_n), .B(n2957), .B(n2957_n), .Y(n3337_n), .Y(n3337) );
 NOR2X1TS U2202 ( .A(n3032), .A(n3032_n), .B(n3216), .B(n3216_n), .Y(n3412_n), .Y(n3412) );
 AND2X2TS U2203 ( .A(n3166), .A(n3166_n), .B(n3422), .B(n3422_n), .Y(n3421_n), .Y(n3421) );
 NOR2X1TS U2204 ( .A(n3423), .A(n3423_n), .B(n3424), .B(n3424_n), .Y(n3422_n), .Y(n3422) );
 NOR2X1TS U2205 ( .A(n3427), .A(n3427_n), .B(n3428), .B(n3428_n), .Y(n3426_n), .Y(n3426) );
 NOR2X1TS U2206 ( .A(n3276), .A(n3276_n), .B(n3432), .B(n3432_n), .Y(n3427_n), .Y(n3427) );
 NOR2X1TS U2207 ( .A(n3433), .A(n3433_n), .B(n3434), .B(n3434_n), .Y(n3425_n), .Y(n3425) );
 NOR2X1TS U2208 ( .A(n3051), .A(n3051_n), .B(n3156), .B(n3156_n), .Y(n3434_n), .Y(n3434) );
 NOR2X1TS U2209 ( .A(n3185), .A(n3185_n), .B(n3435), .B(n3435_n), .Y(n3433_n), .Y(n3433) );
 NOR2X1TS U2210 ( .A(n3439), .A(n3439_n), .B(n3440), .B(n3440_n), .Y(n3436_n), .Y(n3436) );
 INVX2TS U2211 ( .A(n3649), .A(n3649_n), .Y(n3418_n), .Y(n3418) );
 NOR2X1TS U2212 ( .A(n3444), .A(n3444_n), .B(n3445), .B(n3445_n), .Y(n3166_n), .Y(n3166) );
 AND2X2TS U2213 ( .A(n3137), .A(n3137_n), .B(n3448), .B(n3448_n), .Y(n3447_n), .Y(n3447) );
 NOR2X1TS U2214 ( .A(n3450), .A(n3450_n), .B(n3451), .B(n3451_n), .Y(n3446_n), .Y(n3446) );
 NOR2X1TS U2215 ( .A(n3456), .A(n3456_n), .B(n3049), .B(n3049_n), .Y(n3450_n), .Y(n3450) );
 NOR2X1TS U2216 ( .A(n2952), .A(n2952_n), .B(n3458), .B(n3458_n), .Y(n3456_n), .Y(n3456) );
 NOR2X1TS U2217 ( .A(n3461), .A(n3461_n), .B(n3462), .B(n3462_n), .Y(n3460_n), .Y(n3460) );
 NOR2X1TS U2218 ( .A(n3463), .A(n3463_n), .B(n3037), .B(n3037_n), .Y(n3462_n), .Y(n3462) );
 NOR2X1TS U2219 ( .A(n3464), .A(n3464_n), .B(n3006), .B(n3006_n), .Y(n3461_n), .Y(n3461) );
 NOR2X1TS U2220 ( .A(n2956), .A(n2956_n), .B(n3022), .B(n3022_n), .Y(n3464_n), .Y(n3464) );
 NOR2X1TS U2221 ( .A(n3385), .A(n3385_n), .B(n3470), .B(n3470_n), .Y(n3420_n), .Y(n3420) );
 AND2X2TS U2222 ( .A(n3473), .A(n3473_n), .B(n3474), .B(n3474_n), .Y(n3472_n), .Y(n3472) );
 NOR2X1TS U2223 ( .A(n3157), .A(n3157_n), .B(n3475), .B(n3475_n), .Y(n3471_n), .Y(n3471) );
 NOR2X1TS U2224 ( .A(n3020), .A(n3020_n), .B(n3345), .B(n3345_n), .Y(n3475_n), .Y(n3475) );
 NOR2X1TS U2225 ( .A(n3037), .A(n3037_n), .B(n3476), .B(n3476_n), .Y(n3157_n), .Y(n3157) );
 NOR2X1TS U2226 ( .A(n3479), .A(n3479_n), .B(n3480), .B(n3480_n), .Y(n3478_n), .Y(n3478) );
 NOR2X1TS U2227 ( .A(n3483), .A(n3483_n), .B(n3484), .B(n3484_n), .Y(n3481_n), .Y(n3481) );
 NOR2X1TS U2228 ( .A(n3048), .A(n3048_n), .B(n3005), .B(n3005_n), .Y(n3484_n), .Y(n3484) );
 NOR2X1TS U2229 ( .A(n3019), .A(n3019_n), .B(n2951), .B(n2951_n), .Y(n3483_n), .Y(n3483) );
 NOR2X1TS U2230 ( .A(n3153), .A(n3153_n), .B(n3487), .B(n3487_n), .Y(n3485_n), .Y(n3485) );
 NOR2X1TS U2231 ( .A(n3051), .A(n3051_n), .B(n3004), .B(n3004_n), .Y(n3487_n), .Y(n3487) );
 NOR2X1TS U2232 ( .A(n3292), .A(n3292_n), .B(n3488), .B(n3488_n), .Y(n3153_n), .Y(n3153) );
 INVX2TS U2233 ( .A(n3247), .A(n3247_n), .Y(n3292_n), .Y(n3292) );
 AND2X2TS U2234 ( .A(n3489), .A(n3489_n), .B(n3490), .B(n3490_n), .Y(n3477_n), .Y(n3477) );
 NOR2X1TS U2235 ( .A(n3491), .A(n3491_n), .B(n3258), .B(n3258_n), .Y(n3490_n), .Y(n3490) );
 NOR2X1TS U2236 ( .A(n3280), .A(n3280_n), .B(n3492), .B(n3492_n), .Y(n3258_n), .Y(n3258) );
 NOR2X1TS U2237 ( .A(n3493), .A(n3493_n), .B(n3494), .B(n3494_n), .Y(n3489_n), .Y(n3489) );
 NOR2X1TS U2238 ( .A(n3498), .A(n3498_n), .B(n3499), .B(n3499_n), .Y(n3495_n), .Y(n3495) );
 NOR2X1TS U2239 ( .A(n3500), .A(n3500_n), .B(n3501), .B(n3501_n), .Y(n3499_n), .Y(n3499) );
 NOR2X1TS U2240 ( .A(n3502), .A(n3502_n), .B(n3009), .B(n3009_n), .Y(n3498_n), .Y(n3498) );
 NOR2X1TS U2241 ( .A(n3812), .A(n3812_n), .B(n3185), .B(n3185_n), .Y(n3493_n), .Y(n3493) );
 NOR2X1TS U2242 ( .A(n3505), .A(n3505_n), .B(n3506), .B(n3506_n), .Y(n3504_n), .Y(n3504) );
 OR2X2TS U2243 ( .A(n3512), .A(n3512_n), .B(n3513), .B(n3513_n), .Y(n3505_n), .Y(n3505) );
 NOR2X1TS U2244 ( .A(n3516), .A(n3516_n), .B(n3517), .B(n3517_n), .Y(n3503_n), .Y(n3503) );
 NOR2X1TS U2245 ( .A(n3520), .A(n3520_n), .B(n3521), .B(n3521_n), .Y(n3519_n), .Y(n3519) );
 NOR2X1TS U2246 ( .A(n3024), .A(n3024_n), .B(n3277), .B(n3277_n), .Y(n3520_n), .Y(n3520) );
 INVX2TS U2247 ( .A(n2990), .A(n2990_n), .Y(n3277_n), .Y(n3277) );
 NOR2X1TS U2248 ( .A(n3524), .A(n3524_n), .B(n3525), .B(n3525_n), .Y(n3518_n), .Y(n3518) );
 NOR2X1TS U2249 ( .A(n3488), .A(n3488_n), .B(n3319), .B(n3319_n), .Y(n3524_n), .Y(n3524) );
 INVX2TS U2250 ( .A(n2997), .A(n2997_n), .Y(n3488_n), .Y(n3488) );
 NOR2X1TS U2251 ( .A(n3529), .A(n3529_n), .B(n3530), .B(n3530_n), .Y(n3377_n), .Y(n3377) );
 NOR2X1TS U2252 ( .A(n3533), .A(n3533_n), .B(n3534), .B(n3534_n), .Y(n3532_n), .Y(n3532) );
 NOR2X1TS U2253 ( .A(n3052), .A(n3052_n), .B(n3535), .B(n3535_n), .Y(n3533_n), .Y(n3533) );
 NOR2X1TS U2254 ( .A(n3536), .A(n3536_n), .B(n3537), .B(n3537_n), .Y(n3531_n), .Y(n3531) );
 INVX2TS U2255 ( .A(n3540), .A(n3540_n), .Y(n3226_n), .Y(n3226) );
 NOR2X1TS U2256 ( .A(n3543), .A(n3543_n), .B(n3544), .B(n3544_n), .Y(n3542_n), .Y(n3542) );
 NOR2X1TS U2257 ( .A(n3551), .A(n3551_n), .B(n3048), .B(n3048_n), .Y(n3543_n), .Y(n3543) );
 NOR2X1TS U2258 ( .A(n3552), .A(n3552_n), .B(n3553), .B(n3553_n), .Y(n3541_n), .Y(n3541) );
 NOR2X1TS U2259 ( .A(n3560), .A(n3560_n), .B(n3561), .B(n3561_n), .Y(n3559_n), .Y(n3559) );
 NOR2X1TS U2260 ( .A(n3564), .A(n3564_n), .B(n3565), .B(n3565_n), .Y(n3562_n), .Y(n3562) );
 NOR2X1TS U2261 ( .A(n3059), .A(n3059_n), .B(n3568), .B(n3568_n), .Y(n3564_n), .Y(n3564) );
 INVX2TS U2262 ( .A(n3336), .A(n3336_n), .Y(n3568_n), .Y(n3568) );
 NOR2X1TS U2263 ( .A(n3123), .A(n3123_n), .B(n3047), .B(n3047_n), .Y(n3336_n), .Y(n3336) );
 INVX2TS U2264 ( .A(n3626), .A(n3626_n), .Y(n3216_n), .Y(n3216) );
 NOR2X1TS U2265 ( .A(n3571), .A(n3571_n), .B(n3572), .B(n3572_n), .Y(n3558_n), .Y(n3558) );
 OR2X2TS U2266 ( .A(n3573), .A(n3573_n), .B(n3574), .B(n3574_n), .Y(n3572_n), .Y(n3572) );
 NOR2X1TS U2267 ( .A(n3576), .A(n3576_n), .B(n3014), .B(n3014_n), .Y(n3573_n), .Y(n3573) );
 NOR2X1TS U2268 ( .A(n3579), .A(n3579_n), .B(n3580), .B(n3580_n), .Y(n3578_n), .Y(n3578) );
 NOR2X1TS U2269 ( .A(n3086), .A(n3086_n), .B(n2953), .B(n2953_n), .Y(n3579_n), .Y(n3579) );
 NOR2X1TS U2270 ( .A(n3229), .A(n3229_n), .B(n3583), .B(n3583_n), .Y(n3577_n), .Y(n3577) );
 NOR2X1TS U2271 ( .A(n3584), .A(n3584_n), .B(n2987), .B(n2987_n), .Y(n3583_n), .Y(n3583) );
 NOR2X1TS U2272 ( .A(n3585), .A(n3585_n), .B(n3246), .B(n3246_n), .Y(n3584_n), .Y(n3584) );
 NOR2X1TS U2273 ( .A(n3347), .A(n3347_n), .B(n3432), .B(n3432_n), .Y(n3229_n), .Y(n3229) );
 INVX2TS U2274 ( .A(n3586), .A(n3586_n), .Y(n3432_n), .Y(n3432) );
 INVX2TS U2275 ( .A(n2966), .A(n2966_n), .Y(n3347_n), .Y(n3347) );
 OR2X2TS U2276 ( .A(n3589), .A(n3589_n), .B(n3590), .B(n3590_n), .Y(n3281_n), .Y(n3281) );
 NOR2X1TS U2277 ( .A(n3593), .A(n3593_n), .B(n3594), .B(n3594_n), .Y(n3592_n), .Y(n3592) );
 NOR2X1TS U2278 ( .A(n3087), .A(n3087_n), .B(n3218), .B(n3218_n), .Y(n3593_n), .Y(n3593) );
 INVX2TS U2279 ( .A(n2983), .A(n2983_n), .Y(n3218_n), .Y(n3218) );
 NOR2X1TS U2280 ( .A(n3598), .A(n3598_n), .B(n3599), .B(n3599_n), .Y(n3591_n), .Y(n3591) );
 NOR2X1TS U2281 ( .A(n3091), .A(n3091_n), .B(n2954), .B(n2954_n), .Y(n3598_n), .Y(n3598) );
 NOR2X1TS U2282 ( .A(n3604), .A(n3604_n), .B(n3605), .B(n3605_n), .Y(n3603_n), .Y(n3603) );
 NOR2X1TS U2283 ( .A(n3606), .A(n3606_n), .B(n3054), .B(n3054_n), .Y(n3605_n), .Y(n3605) );
 NOR2X1TS U2284 ( .A(n3607), .A(n3607_n), .B(n3024), .B(n3024_n), .Y(n3604_n), .Y(n3604) );
 NOR2X1TS U2285 ( .A(n3376), .A(n3376_n), .B(n3608), .B(n3608_n), .Y(n3607_n), .Y(n3607) );
 INVX2TS U2286 ( .A(n3013), .A(n3013_n), .Y(n3376_n), .Y(n3376) );
 NOR2X1TS U2287 ( .A(n3609), .A(n3609_n), .B(n3610), .B(n3610_n), .Y(n3602_n), .Y(n3602) );
 NOR2X1TS U2288 ( .A(n3613), .A(n3613_n), .B(n3614), .B(n3614_n), .Y(n3611_n), .Y(n3611) );
 NOR2X1TS U2289 ( .A(n2936), .A(n2936_n), .B(n3156), .B(n3156_n), .Y(n3614_n), .Y(n3614) );
 NOR2X1TS U2290 ( .A(n3615), .A(n3615_n), .B(n3050), .B(n3050_n), .Y(n3613_n), .Y(n3613) );
 NOR2X1TS U2291 ( .A(n3266), .A(n3266_n), .B(n3618), .B(n3618_n), .Y(n3617_n), .Y(n3617) );
 AND2X2TS U2292 ( .A(n3268), .A(n3268_n), .B(n3749), .B(n3749_n), .Y(n3620_n), .Y(n3620) );
 NOR2X1TS U2293 ( .A(n3750), .A(n3750_n), .B(n3751), .B(n3751_n), .Y(n3749_n), .Y(n3749) );
 NOR2X1TS U2294 ( .A(n3754), .A(n3754_n), .B(n3755), .B(n3755_n), .Y(n3753_n), .Y(n3753) );
 NOR2X1TS U2295 ( .A(n3368), .A(n3368_n), .B(n2937), .B(n2937_n), .Y(n3755_n), .Y(n3755) );
 NOR2X1TS U2296 ( .A(n2990), .A(n2990_n), .B(n3585), .B(n3585_n), .Y(n3368_n), .Y(n3368) );
 NOR2X1TS U2297 ( .A(n3756), .A(n3756_n), .B(n3085), .B(n3085_n), .Y(n3754_n), .Y(n3754) );
 AND2X2TS U2298 ( .A(n3757), .A(n3757_n), .B(n3468), .B(n3468_n), .Y(n3752_n), .Y(n3752) );
 INVX2TS U2299 ( .A(n3758), .A(n3758_n), .Y(n3373_n), .Y(n3373) );
 NOR2X1TS U2300 ( .A(n3536), .A(n3536_n), .B(n3761), .B(n3761_n), .Y(n3760_n), .Y(n3760) );
 INVX2TS U2301 ( .A(n2960), .A(n2960_n), .Y(n3246_n), .Y(n3246) );
 NOR2X1TS U2302 ( .A(n3053), .A(n3053_n), .B(n2946), .B(n2946_n), .Y(n3536_n), .Y(n3536) );
 NOR2X1TS U2303 ( .A(n3765), .A(n3765_n), .B(n3766), .B(n3766_n), .Y(n3759_n), .Y(n3759) );
 AND2X2TS U2304 ( .A(n3382), .A(n3382_n), .B(n3414), .B(n3414_n), .Y(n3767_n), .Y(n3767) );
 OR2X2TS U2305 ( .A(n3330), .A(n3330_n), .B(n3769), .B(n3769_n), .Y(n3765_n), .Y(n3765) );
 NOR2X1TS U2306 ( .A(n2962), .A(n2962_n), .B(n3719), .B(n3719_n), .Y(n3330_n), .Y(n3330) );
 NOR2X1TS U2307 ( .A(n3770), .A(n3770_n), .B(n3771), .B(n3771_n), .Y(n3268_n), .Y(n3268) );
 NOR2X1TS U2308 ( .A(n3774), .A(n3774_n), .B(n3587), .B(n3587_n), .Y(n3773_n), .Y(n3773) );
 NOR2X1TS U2309 ( .A(n3155), .A(n3155_n), .B(n3768), .B(n3768_n), .Y(n3587_n), .Y(n3587) );
 NOR2X1TS U2310 ( .A(n3738), .A(n3738_n), .B(n3038), .B(n3038_n), .Y(n3774_n), .Y(n3774) );
 INVX2TS U2311 ( .A(n3402), .A(n3402_n), .Y(n3738_n), .Y(n3738) );
 NOR2X1TS U2312 ( .A(n3095), .A(n3095_n), .B(n3540), .B(n3540_n), .Y(n3402_n), .Y(n3402) );
 NOR2X1TS U2313 ( .A(n3775), .A(n3775_n), .B(n3776), .B(n3776_n), .Y(n3772_n), .Y(n3772) );
 NOR2X1TS U2314 ( .A(n3055), .A(n3055_n), .B(n3476), .B(n3476_n), .Y(n3775_n), .Y(n3775) );
 NOR2X1TS U2315 ( .A(n3435), .A(n3435_n), .B(n3719), .B(n3719_n), .Y(n3361_n), .Y(n3361) );
 NOR2X1TS U2316 ( .A(n3780), .A(n3780_n), .B(n3781), .B(n3781_n), .Y(n3778_n), .Y(n3778) );
 AND2X2TS U2317 ( .A(n3352), .A(n3352_n), .B(n3429), .B(n3429_n), .Y(n3788_n), .Y(n3788) );
 NOR2X1TS U2318 ( .A(n3621), .A(n3621_n), .B(n3622), .B(n3622_n), .Y(n3619_n), .Y(n3619) );
 NOR2X1TS U2319 ( .A(n3534), .A(n3534_n), .B(n3625), .B(n3625_n), .Y(n3624_n), .Y(n3624) );
 NOR2X1TS U2320 ( .A(n3016), .A(n3016_n), .B(n3626), .B(n3626_n), .Y(n3625_n), .Y(n3625) );
 NOR2X1TS U2321 ( .A(n3085), .A(n3085_n), .B(n3476), .B(n3476_n), .Y(n3534_n), .Y(n3534) );
 NOR2X1TS U2322 ( .A(n3627), .A(n3627_n), .B(n3628), .B(n3628_n), .Y(n3623_n), .Y(n3623) );
 NOR2X1TS U2323 ( .A(n2986), .A(n2986_n), .B(n3501), .B(n3501_n), .Y(n3628_n), .Y(n3628) );
 NOR2X1TS U2324 ( .A(n3059), .A(n3059_n), .B(n3345), .B(n3345_n), .Y(n3627_n), .Y(n3627) );
 AND2X2TS U2325 ( .A(n3631), .A(n3631_n), .B(n3632), .B(n3632_n), .Y(n3630_n), .Y(n3630) );
 NOR2X1TS U2326 ( .A(n3512), .A(n3512_n), .B(n3633), .B(n3633_n), .Y(n3629_n), .Y(n3629) );
 NOR2X1TS U2327 ( .A(n3634), .A(n3634_n), .B(n3635), .B(n3635_n), .Y(n3633_n), .Y(n3633) );
 NOR2X1TS U2328 ( .A(n2981), .A(n2981_n), .B(n3492), .B(n3492_n), .Y(n3512_n), .Y(n3512) );
 INVX2TS U2329 ( .A(n3550), .A(n3550_n), .Y(n3727_n), .Y(n3727) );
 NOR2X1TS U2330 ( .A(n3638), .A(n3638_n), .B(n3639), .B(n3639_n), .Y(n3637_n), .Y(n3637) );
 NOR2X1TS U2331 ( .A(n3642), .A(n3642_n), .B(n3643), .B(n3643_n), .Y(n3641_n), .Y(n3641) );
 NOR2X1TS U2332 ( .A(n3113), .A(n3113_n), .B(n3118), .B(n3118_n), .Y(n3722_n), .Y(n3722) );
 NOR2X1TS U2333 ( .A(n3647), .A(n3647_n), .B(n3648), .B(n3648_n), .Y(n3644_n), .Y(n3644) );
 NOR2X1TS U2334 ( .A(n3501), .A(n3501_n), .B(n3635), .B(n3635_n), .Y(n3648_n), .Y(n3648) );
 INVX2TS U2335 ( .A(n3067), .A(n3067_n), .Y(n3635_n), .Y(n3635) );
 INVX2TS U2336 ( .A(n2988), .A(n2988_n), .Y(n3501_n), .Y(n3501) );
 NOR2X1TS U2337 ( .A(n3649), .A(n3649_n), .B(n3306), .B(n3306_n), .Y(n3647_n), .Y(n3647) );
 INVX2TS U2338 ( .A(n3042), .A(n3042_n), .Y(n3306_n), .Y(n3306) );
 NOR2X1TS U2339 ( .A(n3082), .A(n3082_n), .B(n2947), .B(n2947_n), .Y(n3649_n), .Y(n3649) );
 NOR2X1TS U2340 ( .A(n3650), .A(n3650_n), .B(n3038), .B(n3038_n), .Y(n3642_n), .Y(n3642) );
 NOR2X1TS U2341 ( .A(n3392), .A(n3392_n), .B(n3301), .B(n3301_n), .Y(n3650_n), .Y(n3650) );
 INVX2TS U2342 ( .A(n2945), .A(n2945_n), .Y(n3301_n), .Y(n3301) );
 INVX2TS U2343 ( .A(n3005), .A(n3005_n), .Y(n3392_n), .Y(n3392) );
 NOR2X1TS U2344 ( .A(n3186), .A(n3186_n), .B(n3651), .B(n3651_n), .Y(n3640_n), .Y(n3640) );
 NOR2X1TS U2345 ( .A(n2970), .A(n2970_n), .B(n3802), .B(n3802_n), .Y(n3653_n), .Y(n3653) );
 AND2X2TS U2346 ( .A(n3342), .A(n3342_n), .B(n3469), .B(n3469_n), .Y(n3652_n), .Y(n3652) );
 NOR2X1TS U2347 ( .A(n3116), .A(n3116_n), .B(n2962), .B(n2962_n), .Y(n3655_n), .Y(n3655) );
 NOR2X1TS U2348 ( .A(n3052), .A(n3052_n), .B(n3095), .B(n3095_n), .Y(n3656_n), .Y(n3656) );
 NOR2X1TS U2349 ( .A(n3657), .A(n3657_n), .B(n3276), .B(n3276_n), .Y(n3186_n), .Y(n3186) );
 NOR2X1TS U2350 ( .A(n3516), .A(n3516_n), .B(n3846), .B(n3846_n), .Y(n3845_n), .Y(n3845) );
 NOR2X1TS U2351 ( .A(n3804), .A(n3804_n), .B(n2970), .B(n2970_n), .Y(n3179_n), .Y(n3179) );
 NOR2X1TS U2352 ( .A(n3122), .A(n3122_n), .B(n3510), .B(n3510_n), .Y(n3233_n), .Y(n3233) );
 NOR2X1TS U2353 ( .A(n2977), .A(n2977_n), .B(n3550), .B(n3550_n), .Y(n3586_n), .Y(n3586) );
 NOR2X1TS U2354 ( .A(n3121), .A(n3121_n), .B(n3757), .B(n3757_n), .Y(n3516_n), .Y(n3516) );
 NOR2X1TS U2355 ( .A(n3407), .A(n3407_n), .B(n3849), .B(n3849_n), .Y(n3844_n), .Y(n3844) );
 NOR2X1TS U2356 ( .A(n3657), .A(n3657_n), .B(n3280), .B(n3280_n), .Y(n3407_n), .Y(n3407) );
 INVX2TS U2357 ( .A(n3348), .A(n3348_n), .Y(n3657_n), .Y(n3657) );
 NOR2X1TS U2358 ( .A(n3549), .A(n3549_n), .B(n3096), .B(n3096_n), .Y(n3348_n), .Y(n3348) );
 AND2X2TS U2359 ( .A(n3658), .A(n3658_n), .B(n3659), .B(n3659_n), .Y(n3636_n), .Y(n3636) );
 NOR2X1TS U2360 ( .A(n3285), .A(n3285_n), .B(n3273), .B(n3273_n), .Y(n3659_n), .Y(n3659) );
 INVX2TS U2361 ( .A(n3476), .A(n3476_n), .Y(n3182_n), .Y(n3182) );
 NOR2X1TS U2362 ( .A(n3664), .A(n3664_n), .B(n3665), .B(n3665_n), .Y(n3658_n), .Y(n3658) );
 INVX2TS U2363 ( .A(n3015), .A(n3015_n), .Y(n3375_n), .Y(n3375) );
 NOR2X1TS U2364 ( .A(n2939), .A(n2939_n), .B(n3049), .B(n3049_n), .Y(n3668_n), .Y(n3668) );
 INVX2TS U2365 ( .A(n3291), .A(n3291_n), .Y(n3419_n), .Y(n3419) );
 NOR2X1TS U2366 ( .A(n3839), .A(n3839_n), .B(n3840), .B(n3840_n), .Y(n3838_n), .Y(n3838) );
 NOR2X1TS U2367 ( .A(n3019), .A(n3019_n), .B(n3013), .B(n3013_n), .Y(n3840_n), .Y(n3840) );
 NOR2X1TS U2368 ( .A(n3454), .A(n3454_n), .B(n3626), .B(n3626_n), .Y(n3839_n), .Y(n3839) );
 NOR2X1TS U2369 ( .A(n2989), .A(n2989_n), .B(n2991), .B(n2991_n), .Y(n3454_n), .Y(n3454) );
 NOR2X1TS U2370 ( .A(n3841), .A(n3841_n), .B(n3842), .B(n3842_n), .Y(n3837_n), .Y(n3837) );
 NOR2X1TS U2371 ( .A(n3058), .A(n3058_n), .B(n3015), .B(n3015_n), .Y(n3841_n), .Y(n3841) );
 NOR2X1TS U2372 ( .A(n3127), .A(n3127_n), .B(n3669), .B(n3669_n), .Y(n3616_n), .Y(n3616) );
 NOR2X1TS U2373 ( .A(n3672), .A(n3672_n), .B(n3673), .B(n3673_n), .Y(n3671_n), .Y(n3671) );
 NOR2X1TS U2374 ( .A(n3793), .A(n3793_n), .B(n3794), .B(n3794_n), .Y(n3670_n), .Y(n3670) );
 NOR2X1TS U2375 ( .A(n3123), .A(n3123_n), .B(n2999), .B(n2999_n), .Y(n3796_n), .Y(n3796) );
 NOR2X1TS U2376 ( .A(n3797), .A(n3797_n), .B(n3798), .B(n3798_n), .Y(n3795_n), .Y(n3795) );
 NOR2X1TS U2377 ( .A(n3802), .A(n3802_n), .B(n2963), .B(n2963_n), .Y(n3257_n), .Y(n3257) );
 NOR2X1TS U2378 ( .A(n3803), .A(n3803_n), .B(n3053), .B(n3053_n), .Y(n3797_n), .Y(n3797) );
 NOR2X1TS U2379 ( .A(n2979), .A(n2979_n), .B(n3001), .B(n3001_n), .Y(n3322_n), .Y(n3322) );
 NOR2X1TS U2380 ( .A(n3113), .A(n3113_n), .B(n3280), .B(n3280_n), .Y(n3597_n), .Y(n3597) );
 INVX2TS U2381 ( .A(n2964), .A(n2964_n), .Y(n3280_n), .Y(n3280) );
 NOR2X1TS U2382 ( .A(n3807), .A(n3807_n), .B(n3491), .B(n3491_n), .Y(n3806_n), .Y(n3806) );
 NOR2X1TS U2383 ( .A(n3057), .A(n3057_n), .B(n3758), .B(n3758_n), .Y(n3491_n), .Y(n3491) );
 NOR2X1TS U2384 ( .A(n3809), .A(n3809_n), .B(n3810), .B(n3810_n), .Y(n3805_n), .Y(n3805) );
 NOR2X1TS U2385 ( .A(n2977), .A(n2977_n), .B(n3091), .B(n3091_n), .Y(n3457_n), .Y(n3457) );
 NOR2X1TS U2386 ( .A(n3297), .A(n3297_n), .B(n3814), .B(n3814_n), .Y(n3813_n), .Y(n3813) );
 NOR2X1TS U2387 ( .A(n3052), .A(n3052_n), .B(n3764), .B(n3764_n), .Y(n3814_n), .Y(n3814) );
 NOR2X1TS U2388 ( .A(n3626), .A(n3626_n), .B(n3035), .B(n3035_n), .Y(n3297_n), .Y(n3297) );
 NOR2X1TS U2389 ( .A(n3678), .A(n3678_n), .B(n3679), .B(n3679_n), .Y(n3677_n), .Y(n3677) );
 INVX2TS U2390 ( .A(n3829), .A(n3829_n), .Y(n3199_n), .Y(n3199) );
 NOR2X1TS U2391 ( .A(n3122), .A(n3122_n), .B(n3549), .B(n3549_n), .Y(n3148_n), .Y(n3148) );
 NOR2X1TS U2392 ( .A(n3681), .A(n3681_n), .B(n3682), .B(n3682_n), .Y(n3680_n), .Y(n3680) );
 INVX2TS U2393 ( .A(n3023), .A(n3023_n), .Y(n3308_n), .Y(n3308) );
 INVX2TS U2394 ( .A(n3812), .A(n3812_n), .Y(n3828_n), .Y(n3828) );
 INVX2TS U2395 ( .A(n3510), .A(n3510_n), .Y(n3465_n), .Y(n3465) );
 INVX2TS U2396 ( .A(n3021), .A(n3021_n), .Y(n3155_n), .Y(n3155) );
 NOR2X1TS U2397 ( .A(n2934), .A(n2934_n), .B(n3271), .B(n3271_n), .Y(n3575_n), .Y(n3575) );
 INVX2TS U2398 ( .A(n3535), .A(n3535_n), .Y(n3271_n), .Y(n3271) );
 NOR2X1TS U2399 ( .A(n3687), .A(n3687_n), .B(n3688), .B(n3688_n), .Y(n3684_n), .Y(n3684) );
 INVX2TS U2400 ( .A(n2933), .A(n2933_n), .Y(n3156_n), .Y(n3156) );
 NOR2X1TS U2401 ( .A(n3691), .A(n3691_n), .B(n3188), .B(n3188_n), .Y(n3689_n), .Y(n3689) );
 NOR2X1TS U2402 ( .A(n3010), .A(n3010_n), .B(n3692), .B(n3692_n), .Y(n3188_n), .Y(n3188) );
 NOR2X1TS U2403 ( .A(n3119), .A(n3119_n), .B(n3029), .B(n3029_n), .Y(n3789_n), .Y(n3789) );
 NOR2X1TS U2404 ( .A(n3500), .A(n3500_n), .B(n3014), .B(n3014_n), .Y(n3691_n), .Y(n3691) );
 NOR2X1TS U2405 ( .A(n3812), .A(n3812_n), .B(n3802), .B(n3802_n), .Y(n3298_n), .Y(n3298) );
 INVX2TS U2406 ( .A(n3785), .A(n3785_n), .Y(n3802_n), .Y(n3802) );
 INVX2TS U2407 ( .A(n2953), .A(n2953_n), .Y(n3449_n), .Y(n3449) );
 NOR2X1TS U2408 ( .A(n3695), .A(n3695_n), .B(n3696), .B(n3696_n), .Y(n3693_n), .Y(n3693) );
 NOR2X1TS U2409 ( .A(n3035), .A(n3035_n), .B(n3049), .B(n3049_n), .Y(n3696_n), .Y(n3696) );
 INVX2TS U2410 ( .A(n3585), .A(n3585_n), .Y(n3345_n), .Y(n3345) );
 NOR2X1TS U2411 ( .A(n3094), .A(n3094_n), .B(n3053), .B(n3053_n), .Y(n3585_n), .Y(n3585) );
 NOR2X1TS U2412 ( .A(n3020), .A(n3020_n), .B(n2960), .B(n2960_n), .Y(n3695_n), .Y(n3695) );
 NOR2X1TS U2413 ( .A(n3697), .A(n3697_n), .B(n3698), .B(n3698_n), .Y(n3204_n), .Y(n3204) );
 NOR2X1TS U2414 ( .A(n3029), .A(n3029_n), .B(n2981), .B(n2981_n), .Y(n3307_n), .Y(n3307) );
 INVX2TS U2415 ( .A(n3147), .A(n3147_n), .Y(n3551_n), .Y(n3551) );
 NOR2X1TS U2416 ( .A(n3702), .A(n3702_n), .B(n3703), .B(n3703_n), .Y(n3699_n), .Y(n3699) );
 NOR2X1TS U2417 ( .A(n3096), .A(n3096_n), .B(n3706), .B(n3706_n), .Y(n3417_n), .Y(n3417) );
 NOR2X1TS U2418 ( .A(n3705), .A(n3705_n), .B(n3311), .B(n3311_n), .Y(n3704_n), .Y(n3704) );
 NOR2X1TS U2419 ( .A(n3706), .A(n3706_n), .B(n3291), .B(n3291_n), .Y(n3311_n), .Y(n3311) );
 INVX2TS U2420 ( .A(n2944), .A(n2944_n), .Y(n3706_n), .Y(n3706) );
 NOR2X1TS U2421 ( .A(n3109), .A(n3109_n), .B(n3869), .B(n3869_n), .Y(n3393_n), .Y(n3393) );
 NOR2X1TS U2422 ( .A(n3014), .A(n3014_n), .B(n3050), .B(n3050_n), .Y(n3705_n), .Y(n3705) );
 NOR2X1TS U2423 ( .A(n3030), .A(n3030_n), .B(n2959), .B(n2959_n), .Y(n3785_n), .Y(n3785) );
 INVX2TS U2424 ( .A(n3054), .A(n3054_n), .Y(n3146_n), .Y(n3146) );
 NOR2X1TS U2425 ( .A(n3053), .A(n3053_n), .B(n2949), .B(n2949_n), .Y(n3702_n), .Y(n3702) );
 NOR2X1TS U2426 ( .A(n2978), .A(n2978_n), .B(n3540), .B(n3540_n), .Y(n3215_n), .Y(n3215) );
 INVX2TS U2427 ( .A(n3784), .A(n3784_n), .Y(n3435_n), .Y(n3435) );
 AND2X2TS U2428 ( .A(n3101), .A(n3101_n), .B(n3099), .B(n3099_n), .Y(n3784_n), .Y(n3784) );
 NOR2X1TS U2429 ( .A(n3709), .A(n3709_n), .B(n3710), .B(n3710_n), .Y(n3708_n), .Y(n3708) );
 INVX2TS U2430 ( .A(n3443), .A(n3443_n), .Y(n3140_n), .Y(n3140) );
 NOR2X1TS U2431 ( .A(n3107), .A(n3107_n), .B(n3105), .B(n3105_n), .Y(n3859_n), .Y(n3859) );
 INVX2TS U2432 ( .A(n3228), .A(n3228_n), .Y(n3372_n), .Y(n3372) );
 NOR2X1TS U2433 ( .A(n3108), .A(n3108_n), .B(n3111), .B(n3111_n), .Y(n3871_n), .Y(n3871) );
 NOR2X1TS U2434 ( .A(n3047), .A(n3047_n), .B(n2945), .B(n2945_n), .Y(n3709_n), .Y(n3709) );
 INVX2TS U2435 ( .A(n3764), .A(n3764_n), .Y(n3198_n), .Y(n3198) );
 NOR2X1TS U2436 ( .A(n3609), .A(n3609_n), .B(n3714), .B(n3714_n), .Y(n3707_n), .Y(n3707) );
 INVX2TS U2437 ( .A(n3858), .A(n3858_n), .Y(n3718_n), .Y(n3718) );
 INVX2TS U2438 ( .A(n3548), .A(n3548_n), .Y(n3713_n), .Y(n3713) );
 NOR2X1TS U2439 ( .A(n3119), .A(n3119_n), .B(n2963), .B(n2963_n), .Y(n3548_n), .Y(n3548) );
 NOR2X1TS U2440 ( .A(n3098), .A(n3098_n), .B(n3102), .B(n3102_n), .Y(n3721_n), .Y(n3721) );
 INVX2TS U2441 ( .A(n3549), .A(n3549_n), .Y(n3654_n), .Y(n3654) );
 NOR2X1TS U2442 ( .A(n3121), .A(n3121_n), .B(n3051), .B(n3051_n), .Y(n3608_n), .Y(n3608) );
 INVX2TS U2443 ( .A(n2994), .A(n2994_n), .Y(n3264_n), .Y(n3264) );
 NOR2X1TS U2444 ( .A(n3104), .A(n3104_n), .B(n3110), .B(n3110_n), .Y(n3877_n), .Y(n3877) );
 NOR2X1TS U2445 ( .A(n3115), .A(n3115_n), .B(n2959), .B(n2959_n), .Y(n3863_n), .Y(n3863) );
 NOR2X1TS U2446 ( .A(n3719), .A(n3719_n), .B(n3720), .B(n3720_n), .Y(n3609_n), .Y(n3609) );
 INVX2TS U2447 ( .A(n3728), .A(n3728_n), .Y(n3719_n), .Y(n3719) );
 NOR2X1TS U2448 ( .A(n2959), .A(n2959_n), .B(n3550), .B(n3550_n), .Y(n3728_n), .Y(n3728) );
 NOR2X1TS U2449 ( .A(n3105), .A(n3105_n), .B(n3106), .B(n3106_n), .Y(n3876_n), .Y(n3876) );
 NAND2BX1TS U2450 ( .AN(n3098), .AN(n3098_n), .B(n3101), .B(n3101_n), .Y(n3812_n), .Y(n3812) );
 NAND2X1TS U2451 ( .A(n3107), .A(n3107_n), .B(n3104), .B(n3104_n), .Y(n3228_n), .Y(n3228) );
 NAND2X1TS U2452 ( .A(n3000), .A(n3000_n), .B(n2959), .B(n2959_n), .Y(n3276_n), .Y(n3276) );
 NOR2BX1TS U2453 ( .AN(n3099), .AN(n3099_n), .B(n3102), .B(n3102_n), .Y(n3184_n), .Y(n3184) );
 NAND2X1TS U2454 ( .A(n3161), .A(n3161_n), .B(n3162), .B(n3162_n), .Y(n3160_n), .Y(n3160) );
 NAND2X1TS U2455 ( .A(n3165), .A(n3165_n), .B(n3166), .B(n3166_n), .Y(n3163_n), .Y(n3163) );
 NAND2X1TS U2456 ( .A(n3169), .A(n3169_n), .B(n3170), .B(n3170_n), .Y(n3168_n), .Y(n3168) );
 NAND2X1TS U2457 ( .A(n3183), .A(n3183_n), .B(n3150), .B(n3150_n), .Y(n3167_n), .Y(n3167) );
 NAND2BX1TS U2458 ( .AN(n3188), .AN(n3188_n), .B(n3189), .B(n3189_n), .Y(n3187_n), .Y(n3187) );
 NAND2X1TS U2459 ( .A(n3190), .A(n3190_n), .B(n3191), .B(n3191_n), .Y(n3159_n), .Y(n3159) );
 NAND2X1TS U2460 ( .A(n3194), .A(n3194_n), .B(n3195), .B(n3195_n), .Y(n3193_n), .Y(n3193) );
 NAND2X1TS U2461 ( .A(n3196), .A(n3196_n), .B(n3197), .B(n3197_n), .Y(n3192_n), .Y(n3192) );
 NAND2X1TS U2462 ( .A(n3043), .A(n3043_n), .B(n2996), .B(n2996_n), .Y(n3197_n), .Y(n3197) );
 NAND2X1TS U2463 ( .A(n3101), .A(n3101_n), .B(n3199), .B(n3199_n), .Y(n3196_n), .Y(n3196) );
 NAND2X1TS U2464 ( .A(n3200), .A(n3200_n), .B(n3201), .B(n3201_n), .Y(d[5]_n), .Y(d[5]) );
 NAND2X1TS U2465 ( .A(n3128), .A(n3128_n), .B(n3204), .B(n3204_n), .Y(n3203_n), .Y(n3203) );
 NAND2X1TS U2466 ( .A(n3236), .A(n3236_n), .B(n3237), .B(n3237_n), .Y(n3202_n), .Y(n3202) );
 NAND2X1TS U2467 ( .A(n3240), .A(n3240_n), .B(n3241), .B(n3241_n), .Y(n3239_n), .Y(n3239) );
 NAND2X1TS U2468 ( .A(n3244), .A(n3244_n), .B(n3245), .B(n3245_n), .Y(n3243_n), .Y(n3243) );
 NAND2X1TS U2469 ( .A(n3081), .A(n3081_n), .B(n2989), .B(n2989_n), .Y(n3245_n), .Y(n3245) );
 NAND2X1TS U2470 ( .A(n2931), .A(n2931_n), .B(n3247), .B(n3247_n), .Y(n3244_n), .Y(n3244) );
 NAND2X1TS U2471 ( .A(n3248), .A(n3248_n), .B(n3249), .B(n3249_n), .Y(n3242_n), .Y(n3242) );
 NAND2X1TS U2472 ( .A(n3066), .A(n3066_n), .B(n3250), .B(n3250_n), .Y(n3249_n), .Y(n3249) );
 NAND2X1TS U2473 ( .A(n2985), .A(n2985_n), .B(n3251), .B(n3251_n), .Y(n3248_n), .Y(n3248) );
 NAND2X1TS U2474 ( .A(n3253), .A(n3253_n), .B(n3254), .B(n3254_n), .Y(n3238_n), .Y(n3238) );
 NAND2X1TS U2475 ( .A(n3146), .A(n3146_n), .B(n3255), .B(n3255_n), .Y(n3254_n), .Y(n3254) );
 NAND2X1TS U2476 ( .A(n3256), .A(n3256_n), .B(n2941), .B(n2941_n), .Y(n3255_n), .Y(n3255) );
 NAND2X1TS U2477 ( .A(n3260), .A(n3260_n), .B(n3261), .B(n3261_n), .Y(n3259_n), .Y(n3259) );
 NAND2X1TS U2478 ( .A(n3075), .A(n3075_n), .B(n3262), .B(n3262_n), .Y(n3261_n), .Y(n3261) );
 NAND2X1TS U2479 ( .A(n3024), .A(n3024_n), .B(n2937), .B(n2937_n), .Y(n3262_n), .Y(n3262) );
 NAND2X1TS U2480 ( .A(n2934), .A(n2934_n), .B(n3263), .B(n3263_n), .Y(n3260_n), .Y(n3260) );
 NAND2X1TS U2481 ( .A(n3264), .A(n3264_n), .B(n3037), .B(n3037_n), .Y(n3263_n), .Y(n3263) );
 NAND2X1TS U2482 ( .A(n3268), .A(n3268_n), .B(n3269), .B(n3269_n), .Y(n3267_n), .Y(n3267) );
 NAND2X1TS U2483 ( .A(n3194), .A(n3194_n), .B(n3731), .B(n3731_n), .Y(n3730_n), .Y(n3730) );
 NAND2X1TS U2484 ( .A(n3486), .A(n3486_n), .B(n3734), .B(n3734_n), .Y(n3733_n), .Y(n3733) );
 NAND2X1TS U2485 ( .A(n3061), .A(n3061_n), .B(n3077), .B(n3077_n), .Y(n3734_n), .Y(n3734) );
 NAND2X1TS U2486 ( .A(n3735), .A(n3735_n), .B(n3736), .B(n3736_n), .Y(n3732_n), .Y(n3732) );
 NAND2X1TS U2487 ( .A(n2932), .A(n2932_n), .B(n2947), .B(n2947_n), .Y(n3736_n), .Y(n3736) );
 NAND2X1TS U2488 ( .A(n3597), .A(n3597_n), .B(n3039), .B(n3039_n), .Y(n3735_n), .Y(n3735) );
 NAND2X1TS U2489 ( .A(n3739), .A(n3739_n), .B(n3740), .B(n3740_n), .Y(n3729_n), .Y(n3729) );
 NAND2X1TS U2490 ( .A(n2990), .A(n2990_n), .B(n3418), .B(n3418_n), .Y(n3742_n), .Y(n3742) );
 NAND2X1TS U2491 ( .A(n3515), .A(n3515_n), .B(n3747), .B(n3747_n), .Y(n3746_n), .Y(n3746) );
 NAND2X1TS U2492 ( .A(n3022), .A(n3022_n), .B(n2942), .B(n2942_n), .Y(n3747_n), .Y(n3747) );
 NAND2X1TS U2493 ( .A(n3051), .A(n3051_n), .B(n3048), .B(n3048_n), .Y(n3272_n), .Y(n3272) );
 NAND2X1TS U2494 ( .A(n3283), .A(n3283_n), .B(n3284), .B(n3284_n), .Y(n3282_n), .Y(n3282) );
 NAND2X1TS U2495 ( .A(n3287), .A(n3287_n), .B(n3288), .B(n3288_n), .Y(n3286_n), .Y(n3286) );
 NAND2X1TS U2496 ( .A(n3008), .A(n3008_n), .B(n3215), .B(n3215_n), .Y(n3288_n), .Y(n3288) );
 NAND2X1TS U2497 ( .A(n3295), .A(n3295_n), .B(n3296), .B(n3296_n), .Y(n3294_n), .Y(n3294) );
 NOR2BX1TS U2498 ( .AN(n3136), .AN(n3136_n), .B(n3297), .B(n3297_n), .Y(n3295_n), .Y(n3295) );
 NAND2X1TS U2499 ( .A(n3299), .A(n3299_n), .B(n3300), .B(n3300_n), .Y(n3293_n), .Y(n3293) );
 NAND2X1TS U2500 ( .A(n3301), .A(n3301_n), .B(n3302), .B(n3302_n), .Y(n3300_n), .Y(n3300) );
 NAND2X1TS U2501 ( .A(n3047), .A(n3047_n), .B(n3089), .B(n3089_n), .Y(n3302_n), .Y(n3302) );
 NAND2X1TS U2502 ( .A(n3124), .A(n3124_n), .B(n3125), .B(n3125_n), .Y(d[7]_n), .Y(d[7]) );
 NAND2X1TS U2503 ( .A(n3128), .A(n3128_n), .B(n3129), .B(n3129_n), .Y(n3126_n), .Y(n3126) );
 NAND2X1TS U2504 ( .A(n3132), .A(n3132_n), .B(n3133), .B(n3133_n), .Y(n3131_n), .Y(n3131) );
 NAND2X1TS U2505 ( .A(n3136), .A(n3136_n), .B(n3137), .B(n3137_n), .Y(n3135_n), .Y(n3135) );
 NAND2X1TS U2506 ( .A(n3044), .A(n3044_n), .B(n3246), .B(n3246_n), .Y(n3136_n), .Y(n3136) );
 NAND2X1TS U2507 ( .A(n3138), .A(n3138_n), .B(n3139), .B(n3139_n), .Y(n3134_n), .Y(n3134) );
 NAND2X1TS U2508 ( .A(n3028), .A(n3028_n), .B(n3140), .B(n3140_n), .Y(n3139_n), .Y(n3139) );
 NAND2X1TS U2509 ( .A(n2969), .A(n2969_n), .B(n3141), .B(n3141_n), .Y(n3138_n), .Y(n3138) );
 NAND2X1TS U2510 ( .A(n3144), .A(n3144_n), .B(n3145), .B(n3145_n), .Y(n3143_n), .Y(n3143) );
 NAND2X1TS U2511 ( .A(n3065), .A(n3065_n), .B(n3147), .B(n3147_n), .Y(n3145_n), .Y(n3145) );
 NAND2X1TS U2512 ( .A(n2964), .A(n2964_n), .B(n3148), .B(n3148_n), .Y(n3144_n), .Y(n3144) );
 NAND2X1TS U2513 ( .A(n3149), .A(n3149_n), .B(n3150), .B(n3150_n), .Y(n3142_n), .Y(n3142) );
 NAND2X1TS U2514 ( .A(n3151), .A(n3151_n), .B(n3152), .B(n3152_n), .Y(n3130_n), .Y(n3130) );
 NAND2X1TS U2515 ( .A(n3207), .A(n3207_n), .B(n3208), .B(n3208_n), .Y(n3206_n), .Y(n3206) );
 NAND2X1TS U2516 ( .A(n3213), .A(n3213_n), .B(n3214), .B(n3214_n), .Y(n3212_n), .Y(n3212) );
 NAND2X1TS U2517 ( .A(n3079), .A(n3079_n), .B(n2950), .B(n2950_n), .Y(n3214_n), .Y(n3214) );
 NAND2X1TS U2518 ( .A(n3070), .A(n3070_n), .B(n3216), .B(n3216_n), .Y(n3213_n), .Y(n3213) );
 NAND2X1TS U2519 ( .A(n3219), .A(n3219_n), .B(n3220), .B(n3220_n), .Y(n3205_n), .Y(n3205) );
 NAND2X1TS U2520 ( .A(n3223), .A(n3223_n), .B(n3224), .B(n3224_n), .Y(n3222_n), .Y(n3222) );
 NAND2X1TS U2521 ( .A(n3067), .A(n3067_n), .B(n3225), .B(n3225_n), .Y(n3224_n), .Y(n3224) );
 NAND2X1TS U2522 ( .A(n3226), .A(n3226_n), .B(n3227), .B(n3227_n), .Y(n3223_n), .Y(n3223) );
 NAND2X1TS U2523 ( .A(n3012), .A(n3012_n), .B(n2940), .B(n2940_n), .Y(n3227_n), .Y(n3227) );
 NAND2X1TS U2524 ( .A(n3231), .A(n3231_n), .B(n3232), .B(n3232_n), .Y(n3230_n), .Y(n3230) );
 NAND2X1TS U2525 ( .A(n3074), .A(n3074_n), .B(n3234), .B(n3234_n), .Y(n3231_n), .Y(n3231) );
 NAND2X1TS U2526 ( .A(n3020), .A(n3020_n), .B(n3235), .B(n3235_n), .Y(n3234_n), .Y(n3234) );
 NAND2X1TS U2527 ( .A(n3792), .A(n3792_n), .B(n3670), .B(n3670_n), .Y(n3791_n), .Y(n3791) );
 NAND2X1TS U2528 ( .A(n3817), .A(n3817_n), .B(n3818), .B(n3818_n), .Y(n3816_n), .Y(n3816) );
 NAND2X1TS U2529 ( .A(n3021), .A(n3021_n), .B(n3819), .B(n3819_n), .Y(n3818_n), .Y(n3818) );
 NAND2X1TS U2530 ( .A(n3256), .A(n3256_n), .B(n3738), .B(n3738_n), .Y(n3819_n), .Y(n3819) );
 NAND2X1TS U2531 ( .A(n3351), .A(n3351_n), .B(n3822), .B(n3822_n), .Y(n3821_n), .Y(n3821) );
 NAND2X1TS U2532 ( .A(n3075), .A(n3075_n), .B(n3823), .B(n3823_n), .Y(n3822_n), .Y(n3822) );
 NAND2X1TS U2533 ( .A(n3826), .A(n3826_n), .B(n3827), .B(n3827_n), .Y(n3815_n), .Y(n3815) );
 NAND2X1TS U2534 ( .A(n3828), .A(n3828_n), .B(n3199), .B(n3199_n), .Y(n3827_n), .Y(n3827) );
 NAND2X1TS U2535 ( .A(n3832), .A(n3832_n), .B(n3833), .B(n3833_n), .Y(n3831_n), .Y(n3831) );
 NAND2X1TS U2536 ( .A(n3017), .A(n3017_n), .B(n3585), .B(n3585_n), .Y(n3833_n), .Y(n3833) );
 NAND2X1TS U2537 ( .A(n3040), .A(n3040_n), .B(n3834), .B(n3834_n), .Y(n3832_n), .Y(n3832) );
 NAND2X1TS U2538 ( .A(n3020), .A(n3020_n), .B(n2986), .B(n2986_n), .Y(n3834_n), .Y(n3834) );
 NAND2X1TS U2539 ( .A(n3473), .A(n3473_n), .B(n3835), .B(n3835_n), .Y(n3830_n), .Y(n3830) );
 NAND2X1TS U2540 ( .A(n2956), .A(n2956_n), .B(n3392), .B(n3392_n), .Y(n3835_n), .Y(n3835) );
 NAND2X1TS U2541 ( .A(n3236), .A(n3236_n), .B(n3836), .B(n3836_n), .Y(n3790_n), .Y(n3790) );
 NAND2X1TS U2542 ( .A(n3854), .A(n3854_n), .B(n3855), .B(n3855_n), .Y(n3853_n), .Y(n3853) );
 NAND2X1TS U2543 ( .A(n3383), .A(n3383_n), .B(n3862), .B(n3862_n), .Y(n3861_n), .Y(n3861) );
 NAND2X1TS U2544 ( .A(n3060), .A(n3060_n), .B(n3021), .B(n3021_n), .Y(n3862_n), .Y(n3862) );
 NAND2X1TS U2545 ( .A(n3864), .A(n3864_n), .B(n3865), .B(n3865_n), .Y(n3852_n), .Y(n3852) );
 NAND2X1TS U2546 ( .A(n3023), .A(n3023_n), .B(n3006), .B(n3006_n), .Y(n3872_n), .Y(n3872) );
 NAND2X1TS U2547 ( .A(n3874), .A(n3874_n), .B(n3875), .B(n3875_n), .Y(n3873_n), .Y(n3873) );
 NAND2X1TS U2548 ( .A(n3017), .A(n3017_n), .B(n3076), .B(n3076_n), .Y(n3875_n), .Y(n3875) );
 NAND2X1TS U2549 ( .A(n3336), .A(n3336_n), .B(n3547), .B(n3547_n), .Y(n3874_n), .Y(n3874) );
 NAND2X1TS U2550 ( .A(n3108), .A(n3108_n), .B(n3085), .B(n3085_n), .Y(n3315_n), .Y(n3315) );
 NAND2X1TS U2551 ( .A(n3319), .A(n3319_n), .B(n3320), .B(n3320_n), .Y(n3318_n), .Y(n3318) );
 NAND2X1TS U2552 ( .A(n3071), .A(n3071_n), .B(n3180), .B(n3180_n), .Y(n3317_n), .Y(n3317) );
 NAND2X1TS U2553 ( .A(n2951), .A(n2951_n), .B(n2940), .B(n2940_n), .Y(n3250_n), .Y(n3250) );
 NAND2X1TS U2554 ( .A(n3325), .A(n3325_n), .B(n3310), .B(n3310_n), .Y(n3324_n), .Y(n3324) );
 NAND2X1TS U2555 ( .A(n3328), .A(n3328_n), .B(n3329), .B(n3329_n), .Y(n3327_n), .Y(n3327) );
 NAND2X1TS U2556 ( .A(n3334), .A(n3334_n), .B(n3335), .B(n3335_n), .Y(n3333_n), .Y(n3333) );
 NAND2X1TS U2557 ( .A(n3082), .A(n3082_n), .B(n3336), .B(n3336_n), .Y(n3335_n), .Y(n3335) );
 NAND2X1TS U2558 ( .A(n3338), .A(n3338_n), .B(n3339), .B(n3339_n), .Y(n3326_n), .Y(n3326) );
 NAND2X1TS U2559 ( .A(n3342), .A(n3342_n), .B(n3343), .B(n3343_n), .Y(n3341_n), .Y(n3341) );
 NAND2X1TS U2560 ( .A(n3066), .A(n3066_n), .B(n3344), .B(n3344_n), .Y(n3343_n), .Y(n3343) );
 NAND2X1TS U2561 ( .A(n2918), .A(n2918_n), .B(n3034), .B(n3034_n), .Y(n3344_n), .Y(n3344) );
 NOR2BX1TS U2562 ( .AN(n3349), .AN(n3349_n), .B(n3350), .B(n3350_n), .Y(n3338_n), .Y(n3338) );
 NAND2X1TS U2563 ( .A(n3351), .A(n3351_n), .B(n3352), .B(n3352_n), .Y(n3350_n), .Y(n3350) );
 NAND2X1TS U2564 ( .A(n3072), .A(n3072_n), .B(n3653), .B(n3653_n), .Y(n3351_n), .Y(n3351) );
 NAND2X1TS U2565 ( .A(n3355), .A(n3355_n), .B(n3356), .B(n3356_n), .Y(n3354_n), .Y(n3354) );
 NAND2X1TS U2566 ( .A(n3094), .A(n3094_n), .B(n3357), .B(n3357_n), .Y(n3356_n), .Y(n3356) );
 NAND2X1TS U2567 ( .A(n3358), .A(n3358_n), .B(n3359), .B(n3359_n), .Y(n3357_n), .Y(n3357) );
 NAND2X1TS U2568 ( .A(n2965), .A(n2965_n), .B(n3360), .B(n3360_n), .Y(n3359_n), .Y(n3359) );
 NAND2X1TS U2569 ( .A(n3718), .A(n3718_n), .B(n3728), .B(n3728_n), .Y(n3355_n), .Y(n3355) );
 NAND2X1TS U2570 ( .A(n3362), .A(n3362_n), .B(n3363), .B(n3363_n), .Y(n3353_n), .Y(n3353) );
 NAND2X1TS U2571 ( .A(n3366), .A(n3366_n), .B(n3367), .B(n3367_n), .Y(n3365_n), .Y(n3365) );
 NAND2X1TS U2572 ( .A(n3072), .A(n3072_n), .B(n2984), .B(n2984_n), .Y(n3367_n), .Y(n3367) );
 NAND2X1TS U2573 ( .A(n2914), .A(n2914_n), .B(n2988), .B(n2988_n), .Y(n3366_n), .Y(n3366) );
 NAND2X1TS U2574 ( .A(n3232), .A(n3232_n), .B(n3371), .B(n3371_n), .Y(n3370_n), .Y(n3370) );
 NAND2X1TS U2575 ( .A(n3060), .A(n3060_n), .B(n3372), .B(n3372_n), .Y(n3371_n), .Y(n3371) );
 NAND2X1TS U2576 ( .A(n3081), .A(n3081_n), .B(n3373), .B(n3373_n), .Y(n3232_n), .Y(n3232) );
 NAND2X1TS U2577 ( .A(n3377), .A(n3377_n), .B(n3378), .B(n3378_n), .Y(n3323_n), .Y(n3323) );
 NAND2X1TS U2578 ( .A(n3381), .A(n3381_n), .B(n3382), .B(n3382_n), .Y(n3380_n), .Y(n3380) );
 NAND2X1TS U2579 ( .A(n3026), .A(n3026_n), .B(n3042), .B(n3042_n), .Y(n3383_n), .Y(n3383) );
 NAND2X1TS U2580 ( .A(n3387), .A(n3387_n), .B(n3388), .B(n3388_n), .Y(n3270_n), .Y(n3270) );
 NAND2X1TS U2581 ( .A(n3391), .A(n3391_n), .B(n3241), .B(n3241_n), .Y(n3390_n), .Y(n3390) );
 NAND2X1TS U2582 ( .A(n3392), .A(n3392_n), .B(n3393), .B(n3393_n), .Y(n3241_n), .Y(n3241) );
 NAND2X1TS U2583 ( .A(n3394), .A(n3394_n), .B(n3395), .B(n3395_n), .Y(n3389_n), .Y(n3389) );
 NAND2X1TS U2584 ( .A(n3146), .A(n3146_n), .B(n3396), .B(n3396_n), .Y(n3395_n), .Y(n3395) );
 NAND2X1TS U2585 ( .A(n3400), .A(n3400_n), .B(n3401), .B(n3401_n), .Y(n3399_n), .Y(n3399) );
 NAND2BX1TS U2586 ( .AN(n3217), .AN(n3217_n), .B(n3402), .B(n3402_n), .Y(n3401_n), .Y(n3401) );
 NAND2X1TS U2587 ( .A(n3376), .A(n3376_n), .B(n3403), .B(n3403_n), .Y(n3400_n), .Y(n3400) );
 NAND2X1TS U2588 ( .A(n3057), .A(n3057_n), .B(n3050), .B(n3050_n), .Y(n3403_n), .Y(n3403) );
 NAND2X1TS U2589 ( .A(n3404), .A(n3404_n), .B(n3405), .B(n3405_n), .Y(n3398_n), .Y(n3398) );
 NAND2X1TS U2590 ( .A(n3078), .A(n3078_n), .B(n3406), .B(n3406_n), .Y(n3405_n), .Y(n3405) );
 NAND2X1TS U2591 ( .A(n2908), .A(n2908_n), .B(n2946), .B(n2946_n), .Y(n3406_n), .Y(n3406) );
 NAND2X1TS U2592 ( .A(n2989), .A(n2989_n), .B(n2948), .B(n2948_n), .Y(n3413_n), .Y(n3413) );
 NAND2X1TS U2593 ( .A(n3040), .A(n3040_n), .B(n3418), .B(n3418_n), .Y(n3416_n), .Y(n3416) );
 NAND2X1TS U2594 ( .A(n3419), .A(n3419_n), .B(n3141), .B(n3141_n), .Y(n3415_n), .Y(n3415) );
 NAND2X1TS U2595 ( .A(n3420), .A(n3420_n), .B(n3421), .B(n3421_n), .Y(n3309_n), .Y(n3309) );
 NAND2X1TS U2596 ( .A(n3425), .A(n3425_n), .B(n3426), .B(n3426_n), .Y(n3424_n), .Y(n3424) );
 NAND2X1TS U2597 ( .A(n3429), .A(n3429_n), .B(n3430), .B(n3430_n), .Y(n3428_n), .Y(n3428) );
 NAND2X1TS U2598 ( .A(n3070), .A(n3070_n), .B(n3431), .B(n3431_n), .Y(n3430_n), .Y(n3430) );
 NAND2X1TS U2599 ( .A(n3058), .A(n3058_n), .B(n3320), .B(n3320_n), .Y(n3431_n), .Y(n3431) );
 NAND2X1TS U2600 ( .A(n3436), .A(n3436_n), .B(n3437), .B(n3437_n), .Y(n3423_n), .Y(n3423) );
 NAND2X1TS U2601 ( .A(n3301), .A(n3301_n), .B(n3438), .B(n3438_n), .Y(n3437_n), .Y(n3437) );
 NAND2X1TS U2602 ( .A(n3441), .A(n3441_n), .B(n3442), .B(n3442_n), .Y(n3440_n), .Y(n3440) );
 NAND2X1TS U2603 ( .A(n3039), .A(n3039_n), .B(n2984), .B(n2984_n), .Y(n3442_n), .Y(n3442) );
 NAND2X1TS U2604 ( .A(n3246), .A(n3246_n), .B(n3418), .B(n3418_n), .Y(n3441_n), .Y(n3441) );
 NAND2X1TS U2605 ( .A(n3446), .A(n3446_n), .B(n3447), .B(n3447_n), .Y(n3445_n), .Y(n3445) );
 NAND2X1TS U2606 ( .A(n3402), .A(n3402_n), .B(n3065), .B(n3065_n), .Y(n3448_n), .Y(n3448) );
 NAND2X1TS U2607 ( .A(n2994), .A(n2994_n), .B(n3449), .B(n3449_n), .Y(n3137_n), .Y(n3137) );
 NAND2X1TS U2608 ( .A(n3452), .A(n3452_n), .B(n3453), .B(n3453_n), .Y(n3451_n), .Y(n3451) );
 NAND2BX1TS U2609 ( .AN(n3454), .AN(n3454_n), .B(n3083), .B(n3083_n), .Y(n3453_n), .Y(n3453) );
 NAND2X1TS U2610 ( .A(n3068), .A(n3068_n), .B(n3455), .B(n3455_n), .Y(n3452_n), .Y(n3452) );
 NAND2X1TS U2611 ( .A(n3012), .A(n3012_n), .B(n3015), .B(n3015_n), .Y(n3455_n), .Y(n3455) );
 NAND2X1TS U2612 ( .A(n3010), .A(n3010_n), .B(n3035), .B(n3035_n), .Y(n3458_n), .Y(n3458) );
 NAND2X1TS U2613 ( .A(n3459), .A(n3459_n), .B(n3460), .B(n3460_n), .Y(n3444_n), .Y(n3444) );
 NOR2BX1TS U2614 ( .AN(n3466), .AN(n3466_n), .B(n3467), .B(n3467_n), .Y(n3459_n), .Y(n3459) );
 NAND2X1TS U2615 ( .A(n3468), .A(n3468_n), .B(n3469), .B(n3469_n), .Y(n3467_n), .Y(n3467) );
 NAND2X1TS U2616 ( .A(n3471), .A(n3471_n), .B(n3472), .B(n3472_n), .Y(n3470_n), .Y(n3470) );
 NAND2X1TS U2617 ( .A(n3336), .A(n3336_n), .B(n2914), .B(n2914_n), .Y(n3474_n), .Y(n3474) );
 NAND2X1TS U2618 ( .A(n3654), .A(n3654_n), .B(n2975), .B(n2975_n), .Y(n3473_n), .Y(n3473) );
 NAND2X1TS U2619 ( .A(n3477), .A(n3477_n), .B(n3478), .B(n3478_n), .Y(n3385_n), .Y(n3385) );
 NAND2X1TS U2620 ( .A(n3481), .A(n3481_n), .B(n3482), .B(n3482_n), .Y(n3480_n), .Y(n3480) );
 NAND2X1TS U2621 ( .A(n3485), .A(n3485_n), .B(n3486), .B(n3486_n), .Y(n3479_n), .Y(n3479) );
 NAND2X1TS U2622 ( .A(n2944), .A(n2944_n), .B(n3182), .B(n3182_n), .Y(n3486_n), .Y(n3486) );
 NAND2X1TS U2623 ( .A(n3059), .A(n3059_n), .B(n3023), .B(n3023_n), .Y(n3247_n), .Y(n3247) );
 NAND2X1TS U2624 ( .A(n3495), .A(n3495_n), .B(n3496), .B(n3496_n), .Y(n3494_n), .Y(n3494) );
 NAND2X1TS U2625 ( .A(n3017), .A(n3017_n), .B(n3497), .B(n3497_n), .Y(n3496_n), .Y(n3496) );
 NAND2X1TS U2626 ( .A(n3013), .A(n3013_n), .B(n3488), .B(n3488_n), .Y(n3497_n), .Y(n3497) );
 NAND2X1TS U2627 ( .A(n3348), .A(n3348_n), .B(n3118), .B(n3118_n), .Y(n3185_n), .Y(n3185) );
 NAND2X1TS U2628 ( .A(n3503), .A(n3503_n), .B(n3504), .B(n3504_n), .Y(n3386_n), .Y(n3386) );
 NAND2X1TS U2629 ( .A(n3507), .A(n3507_n), .B(n3508), .B(n3508_n), .Y(n3506_n), .Y(n3506) );
 NAND2X1TS U2630 ( .A(n3298), .A(n3298_n), .B(n3509), .B(n3509_n), .Y(n3508_n), .Y(n3508) );
 NAND2X1TS U2631 ( .A(n3510), .A(n3510_n), .B(n3345), .B(n3345_n), .Y(n3509_n), .Y(n3509) );
 NAND2X1TS U2632 ( .A(n3065), .A(n3065_n), .B(n3511), .B(n3511_n), .Y(n3507_n), .Y(n3507) );
 NAND2X1TS U2633 ( .A(n2949), .A(n2949_n), .B(n3149), .B(n3149_n), .Y(n3511_n), .Y(n3511) );
 NAND2X1TS U2634 ( .A(n2993), .A(n2993_n), .B(n2976), .B(n2976_n), .Y(n3149_n), .Y(n3149) );
 NAND2X1TS U2635 ( .A(n3514), .A(n3514_n), .B(n3515), .B(n3515_n), .Y(n3513_n), .Y(n3513) );
 NAND2X1TS U2636 ( .A(n3026), .A(n3026_n), .B(n3608), .B(n3608_n), .Y(n3515_n), .Y(n3515) );
 NAND2X1TS U2637 ( .A(n3518), .A(n3518_n), .B(n3519), .B(n3519_n), .Y(n3517_n), .Y(n3517) );
 NAND2X1TS U2638 ( .A(n3522), .A(n3522_n), .B(n3523), .B(n3523_n), .Y(n3521_n), .Y(n3521) );
 NAND2X1TS U2639 ( .A(n3027), .A(n3027_n), .B(n2933), .B(n2933_n), .Y(n3523_n), .Y(n3523) );
 NAND2X1TS U2640 ( .A(n3025), .A(n3025_n), .B(n3417), .B(n3417_n), .Y(n3522_n), .Y(n3522) );
 NAND2X1TS U2641 ( .A(n3526), .A(n3526_n), .B(n3527), .B(n3527_n), .Y(n3525_n), .Y(n3525) );
 NAND2X1TS U2642 ( .A(n3081), .A(n3081_n), .B(n3528), .B(n3528_n), .Y(n3527_n), .Y(n3527) );
 NAND2X1TS U2643 ( .A(n3070), .A(n3070_n), .B(n3179), .B(n3179_n), .Y(n3526_n), .Y(n3526) );
 NAND2X1TS U2644 ( .A(n3531), .A(n3531_n), .B(n3532), .B(n3532_n), .Y(n3530_n), .Y(n3530) );
 NAND2X1TS U2645 ( .A(n3538), .A(n3538_n), .B(n3539), .B(n3539_n), .Y(n3537_n), .Y(n3537) );
 NAND2X1TS U2646 ( .A(n3226), .A(n3226_n), .B(n3043), .B(n3043_n), .Y(n3539_n), .Y(n3539) );
 NAND2X1TS U2647 ( .A(n2991), .A(n2991_n), .B(n3067), .B(n3067_n), .Y(n3538_n), .Y(n3538) );
 NAND2X1TS U2648 ( .A(n3541), .A(n3541_n), .B(n3542), .B(n3542_n), .Y(n3529_n), .Y(n3529) );
 NAND2X1TS U2649 ( .A(n3545), .A(n3545_n), .B(n3546), .B(n3546_n), .Y(n3544_n), .Y(n3544) );
 NAND2X1TS U2650 ( .A(n2932), .A(n2932_n), .B(n3547), .B(n3547_n), .Y(n3546_n), .Y(n3546) );
 NAND2X1TS U2651 ( .A(n3019), .A(n3019_n), .B(n3058), .B(n3058_n), .Y(n3547_n), .Y(n3547) );
 NAND2X1TS U2652 ( .A(n3548), .A(n3548_n), .B(n3360), .B(n3360_n), .Y(n3545_n), .Y(n3545) );
 NAND2X1TS U2653 ( .A(n3549), .A(n3549_n), .B(n3550), .B(n3550_n), .Y(n3360_n), .Y(n3360) );
 NAND2X1TS U2654 ( .A(n3554), .A(n3554_n), .B(n3555), .B(n3555_n), .Y(n3553_n), .Y(n3553) );
 NAND2X1TS U2655 ( .A(n3032), .A(n3032_n), .B(n3556), .B(n3556_n), .Y(n3555_n), .Y(n3555) );
 NAND2X1TS U2656 ( .A(n3009), .A(n3009_n), .B(n2961), .B(n2961_n), .Y(n3556_n), .Y(n3556) );
 NAND2X1TS U2657 ( .A(n3558), .A(n3558_n), .B(n3559), .B(n3559_n), .Y(n3164_n), .Y(n3164) );
 NAND2X1TS U2658 ( .A(n3562), .A(n3562_n), .B(n3563), .B(n3563_n), .Y(n3561_n), .Y(n3561) );
 NAND2X1TS U2659 ( .A(n3064), .A(n3064_n), .B(n2983), .B(n2983_n), .Y(n3563_n), .Y(n3563) );
 NAND2X1TS U2660 ( .A(n3566), .A(n3566_n), .B(n3567), .B(n3567_n), .Y(n3565_n), .Y(n3565) );
 NAND2X1TS U2661 ( .A(n3569), .A(n3569_n), .B(n3570), .B(n3570_n), .Y(n3560_n), .Y(n3560) );
 NAND2X1TS U2662 ( .A(n3028), .A(n3028_n), .B(n3060), .B(n3060_n), .Y(n3570_n), .Y(n3570) );
 NAND2X1TS U2663 ( .A(n2993), .A(n2993_n), .B(n2998), .B(n2998_n), .Y(n3569_n), .Y(n3569) );
 NAND2X1TS U2664 ( .A(n3577), .A(n3577_n), .B(n3578), .B(n3578_n), .Y(n3571_n), .Y(n3571) );
 NAND2X1TS U2665 ( .A(n3581), .A(n3581_n), .B(n3582), .B(n3582_n), .Y(n3580_n), .Y(n3580) );
 NAND2X1TS U2666 ( .A(n3042), .A(n3042_n), .B(n2985), .B(n2985_n), .Y(n3582_n), .Y(n3582) );
 NAND2X1TS U2667 ( .A(n3072), .A(n3072_n), .B(n3198), .B(n3198_n), .Y(n3581_n), .Y(n3581) );
 NAND2X1TS U2668 ( .A(n3591), .A(n3591_n), .B(n3592), .B(n3592_n), .Y(n3590_n), .Y(n3590) );
 NAND2X1TS U2669 ( .A(n3595), .A(n3595_n), .B(n3596), .B(n3596_n), .Y(n3594_n), .Y(n3594) );
 NAND2X1TS U2670 ( .A(n3076), .A(n3076_n), .B(n3597), .B(n3597_n), .Y(n3596_n), .Y(n3596) );
 NAND2X1TS U2671 ( .A(n3600), .A(n3600_n), .B(n3601), .B(n3601_n), .Y(n3599_n), .Y(n3599) );
 NAND2X1TS U2672 ( .A(n3067), .A(n3067_n), .B(n3246), .B(n3246_n), .Y(n3600_n), .Y(n3600) );
 NAND2X1TS U2673 ( .A(n3602), .A(n3602_n), .B(n3603), .B(n3603_n), .Y(n3589_n), .Y(n3589) );
 NAND2X1TS U2674 ( .A(n3611), .A(n3611_n), .B(n3612), .B(n3612_n), .Y(n3610_n), .Y(n3610) );
 NAND2X1TS U2675 ( .A(n2994), .A(n2994_n), .B(n2973), .B(n2973_n), .Y(n3612_n), .Y(n3612) );
 NAND2X1TS U2676 ( .A(n3616), .A(n3616_n), .B(n3617), .B(n3617_n), .Y(d[1]_n), .Y(d[1]) );
 NAND2X1TS U2677 ( .A(n3619), .A(n3619_n), .B(n3620), .B(n3620_n), .Y(n3618_n), .Y(n3618) );
 NAND2X1TS U2678 ( .A(n3752), .A(n3752_n), .B(n3753), .B(n3753_n), .Y(n3751_n), .Y(n3751) );
 NAND2X1TS U2679 ( .A(n3032), .A(n3032_n), .B(n3373), .B(n3373_n), .Y(n3468_n), .Y(n3468) );
 NAND2X1TS U2680 ( .A(n3759), .A(n3759_n), .B(n3760), .B(n3760_n), .Y(n3750_n), .Y(n3750) );
 NAND2X1TS U2681 ( .A(n3762), .A(n3762_n), .B(n3763), .B(n3763_n), .Y(n3761_n), .Y(n3761) );
 NAND2X1TS U2682 ( .A(n2931), .A(n2931_n), .B(n2947), .B(n2947_n), .Y(n3763_n), .Y(n3763) );
 NAND2X1TS U2683 ( .A(n3018), .A(n3018_n), .B(n3225), .B(n3225_n), .Y(n3762_n), .Y(n3762) );
 NAND2X1TS U2684 ( .A(n3016), .A(n3016_n), .B(n2960), .B(n2960_n), .Y(n3225_n), .Y(n3225) );
 NAND2X1TS U2685 ( .A(n3767), .A(n3767_n), .B(n3482), .B(n3482_n), .Y(n3766_n), .Y(n3766) );
 NAND2X1TS U2686 ( .A(n3079), .A(n3079_n), .B(n2968), .B(n2968_n), .Y(n3482_n), .Y(n3482) );
 NAND2X1TS U2687 ( .A(n3072), .A(n3072_n), .B(n3002), .B(n3002_n), .Y(n3414_n), .Y(n3414) );
 NAND2X1TS U2688 ( .A(n3041), .A(n3041_n), .B(n3068), .B(n3068_n), .Y(n3382_n), .Y(n3382) );
 NAND2X1TS U2689 ( .A(n3195), .A(n3195_n), .B(n3384), .B(n3384_n), .Y(n3769_n), .Y(n3769) );
 NAND2X1TS U2690 ( .A(n2975), .A(n2975_n), .B(n3727), .B(n3727_n), .Y(n3384_n), .Y(n3384) );
 NAND2X1TS U2691 ( .A(n2995), .A(n2995_n), .B(n3061), .B(n3061_n), .Y(n3195_n), .Y(n3195) );
 NAND2X1TS U2692 ( .A(n3772), .A(n3772_n), .B(n3773), .B(n3773_n), .Y(n3771_n), .Y(n3771) );
 NAND2X1TS U2693 ( .A(n3601), .A(n3601_n), .B(n3777), .B(n3777_n), .Y(n3776_n), .Y(n3776) );
 NAND2X1TS U2694 ( .A(n3375), .A(n3375_n), .B(n3045), .B(n3045_n), .Y(n3777_n), .Y(n3777) );
 NAND2X1TS U2695 ( .A(n3026), .A(n3026_n), .B(n2988), .B(n2988_n), .Y(n3601_n), .Y(n3601) );
 NAND2X1TS U2696 ( .A(n3778), .A(n3778_n), .B(n3779), .B(n3779_n), .Y(n3770_n), .Y(n3770) );
 NAND2X1TS U2697 ( .A(n3123), .A(n3123_n), .B(n3361), .B(n3361_n), .Y(n3779_n), .Y(n3779) );
 NAND2X1TS U2698 ( .A(n3782), .A(n3782_n), .B(n3783), .B(n3783_n), .Y(n3781_n), .Y(n3781) );
 NAND2X1TS U2699 ( .A(n2948), .A(n2948_n), .B(n3528), .B(n3528_n), .Y(n3783_n), .Y(n3783) );
 NAND2X1TS U2700 ( .A(n3011), .A(n3011_n), .B(n3009), .B(n3009_n), .Y(n3528_n), .Y(n3528) );
 NAND2X1TS U2701 ( .A(n3071), .A(n3071_n), .B(n3786), .B(n3786_n), .Y(n3782_n), .Y(n3782) );
 NAND2X1TS U2702 ( .A(n3787), .A(n3787_n), .B(n3764), .B(n3764_n), .Y(n3786_n), .Y(n3786) );
 NAND2X1TS U2703 ( .A(n3788), .A(n3788_n), .B(n3554), .B(n3554_n), .Y(n3780_n), .Y(n3780) );
 NAND2X1TS U2704 ( .A(n2980), .A(n2980_n), .B(n3148), .B(n3148_n), .Y(n3554_n), .Y(n3554) );
 NAND2X1TS U2705 ( .A(n3083), .A(n3083_n), .B(n3656), .B(n3656_n), .Y(n3429_n), .Y(n3429) );
 NAND2BX1TS U2706 ( .AN(n3692), .AN(n3692_n), .B(n3076), .B(n3076_n), .Y(n3352_n), .Y(n3352) );
 NAND2X1TS U2707 ( .A(n3623), .A(n3623_n), .B(n3624), .B(n3624_n), .Y(n3622_n), .Y(n3622) );
 NAND2X1TS U2708 ( .A(n3629), .A(n3629_n), .B(n3630), .B(n3630_n), .Y(n3621_n), .Y(n3621) );
 NAND2X1TS U2709 ( .A(n3021), .A(n3021_n), .B(n2957), .B(n2957_n), .Y(n3632_n), .Y(n3632) );
 NAND2X1TS U2710 ( .A(n3045), .A(n3045_n), .B(n3314), .B(n3314_n), .Y(n3631_n), .Y(n3631) );
 NAND2X1TS U2711 ( .A(n3501), .A(n3501_n), .B(n2939), .B(n2939_n), .Y(n3314_n), .Y(n3314) );
 NAND2X1TS U2712 ( .A(n2977), .A(n2977_n), .B(n3727), .B(n3727_n), .Y(n3492_n), .Y(n3492) );
 NAND2X1TS U2713 ( .A(n3636), .A(n3636_n), .B(n3637), .B(n3637_n), .Y(n3266_n), .Y(n3266) );
 NAND2X1TS U2714 ( .A(n3640), .A(n3640_n), .B(n3641), .B(n3641_n), .Y(n3639_n), .Y(n3639) );
 NAND2X1TS U2715 ( .A(n3644), .A(n3644_n), .B(n3645), .B(n3645_n), .Y(n3643_n), .Y(n3643) );
 NAND2X1TS U2716 ( .A(n3070), .A(n3070_n), .B(n3646), .B(n3646_n), .Y(n3645_n), .Y(n3645) );
 NAND2X1TS U2717 ( .A(n3540), .A(n3540_n), .B(n3320), .B(n3320_n), .Y(n3646_n), .Y(n3646) );
 NAND2X1TS U2718 ( .A(n3721), .A(n3721_n), .B(n3722), .B(n3722_n), .Y(n3320_n), .Y(n3320) );
 NAND2X1TS U2719 ( .A(n3652), .A(n3652_n), .B(n3514), .B(n3514_n), .Y(n3651_n), .Y(n3651) );
 NAND2X1TS U2720 ( .A(n3075), .A(n3075_n), .B(n3653), .B(n3653_n), .Y(n3514_n), .Y(n3514) );
 NAND2X1TS U2721 ( .A(n3654), .A(n3654_n), .B(n3655), .B(n3655_n), .Y(n3469_n), .Y(n3469) );
 NAND2X1TS U2722 ( .A(n3026), .A(n3026_n), .B(n3656), .B(n3656_n), .Y(n3342_n), .Y(n3342) );
 NAND2X1TS U2723 ( .A(n3844), .A(n3844_n), .B(n3845), .B(n3845_n), .Y(n3638_n), .Y(n3638) );
 NAND2X1TS U2724 ( .A(n3847), .A(n3847_n), .B(n3848), .B(n3848_n), .Y(n3846_n), .Y(n3846) );
 NAND2X1TS U2725 ( .A(n3074), .A(n3074_n), .B(n3179), .B(n3179_n), .Y(n3848_n), .Y(n3848) );
 NAND2X1TS U2726 ( .A(n3586), .A(n3586_n), .B(n3824), .B(n3824_n), .Y(n3847_n), .Y(n3847) );
 NOR2BX1TS U2727 ( .AN(n3098), .AN(n3098_n), .B(n3117), .B(n3117_n), .Y(n3824_n), .Y(n3824) );
 NAND2X1TS U2728 ( .A(n3828), .A(n3828_n), .B(n3728), .B(n3728_n), .Y(n3757_n), .Y(n3757) );
 NAND2X1TS U2729 ( .A(n3466), .A(n3466_n), .B(n3850), .B(n3850_n), .Y(n3849_n), .Y(n3849) );
 NAND2X1TS U2730 ( .A(n3438), .A(n3438_n), .B(n3851), .B(n3851_n), .Y(n3850_n), .Y(n3850) );
 NAND2X1TS U2731 ( .A(n3005), .A(n3005_n), .B(n3004), .B(n3004_n), .Y(n3851_n), .Y(n3851) );
 NAND2X1TS U2732 ( .A(n3052), .A(n3052_n), .B(n3087), .B(n3087_n), .Y(n3438_n), .Y(n3438) );
 NAND2X1TS U2733 ( .A(n3148), .A(n3148_n), .B(n2967), .B(n2967_n), .Y(n3466_n), .Y(n3466) );
 NAND2X1TS U2734 ( .A(n3660), .A(n3660_n), .B(n3661), .B(n3661_n), .Y(n3273_n), .Y(n3273) );
 NAND2X1TS U2735 ( .A(n3041), .A(n3041_n), .B(n3002), .B(n3002_n), .Y(n3661_n), .Y(n3661) );
 NAND2X1TS U2736 ( .A(n3465), .A(n3465_n), .B(n3182), .B(n3182_n), .Y(n3660_n), .Y(n3660) );
 NAND2X1TS U2737 ( .A(n3114), .A(n3114_n), .B(n2974), .B(n2974_n), .Y(n3476_n), .Y(n3476) );
 NAND2X1TS U2738 ( .A(n3662), .A(n3662_n), .B(n3663), .B(n3663_n), .Y(n3285_n), .Y(n3285) );
 NAND2X1TS U2739 ( .A(n3077), .A(n3077_n), .B(n3449), .B(n3449_n), .Y(n3663_n), .Y(n3663) );
 NAND2X1TS U2740 ( .A(n3007), .A(n3007_n), .B(n3271), .B(n3271_n), .Y(n3662_n), .Y(n3662) );
 NAND2X1TS U2741 ( .A(n3666), .A(n3666_n), .B(n3667), .B(n3667_n), .Y(n3665_n), .Y(n3665) );
 NAND2X1TS U2742 ( .A(n3082), .A(n3082_n), .B(n3375), .B(n3375_n), .Y(n3667_n), .Y(n3667) );
 NOR2BX1TS U2743 ( .AN(n3567), .AN(n3567_n), .B(n3668), .B(n3668_n), .Y(n3666_n), .Y(n3666) );
 NAND2X1TS U2744 ( .A(n2956), .A(n2956_n), .B(n3419), .B(n3419_n), .Y(n3567_n), .Y(n3567) );
 NAND2X1TS U2745 ( .A(n3837), .A(n3837_n), .B(n3838), .B(n3838_n), .Y(n3664_n), .Y(n3664) );
 NAND2X1TS U2746 ( .A(n3588), .A(n3588_n), .B(n3843), .B(n3843_n), .Y(n3842_n), .Y(n3842) );
 NAND2X1TS U2747 ( .A(n3064), .A(n3064_n), .B(n3062), .B(n3062_n), .Y(n3843_n), .Y(n3843) );
 NAND2X1TS U2748 ( .A(n3308), .A(n3308_n), .B(n2952), .B(n2952_n), .Y(n3588_n), .Y(n3588) );
 NAND2X1TS U2749 ( .A(n3670), .A(n3670_n), .B(n3671), .B(n3671_n), .Y(n3669_n), .Y(n3669) );
 NAND2X1TS U2750 ( .A(n3566), .A(n3566_n), .B(n3674), .B(n3674_n), .Y(n3673_n), .Y(n3673) );
 NAND2X1TS U2751 ( .A(n3027), .A(n3027_n), .B(n2968), .B(n2968_n), .Y(n3674_n), .Y(n3674) );
 NAND2X1TS U2752 ( .A(n3002), .A(n3002_n), .B(n3095), .B(n3095_n), .Y(n3768_n), .Y(n3768) );
 NAND2X1TS U2753 ( .A(n2995), .A(n2995_n), .B(n3308), .B(n3308_n), .Y(n3566_n), .Y(n3566) );
 NAND2X1TS U2754 ( .A(n3675), .A(n3675_n), .B(n3676), .B(n3676_n), .Y(n3672_n), .Y(n3672) );
 NAND2X1TS U2755 ( .A(n2967), .A(n2967_n), .B(n3039), .B(n3039_n), .Y(n3676_n), .Y(n3676) );
 NAND2X1TS U2756 ( .A(n3079), .A(n3079_n), .B(n3003), .B(n3003_n), .Y(n3675_n), .Y(n3675) );
 NAND2X1TS U2757 ( .A(n3548), .A(n3548_n), .B(n3029), .B(n3029_n), .Y(n3174_n), .Y(n3174) );
 NAND2X1TS U2758 ( .A(n3795), .A(n3795_n), .B(n3349), .B(n3349_n), .Y(n3794_n), .Y(n3794) );
 NAND2X1TS U2759 ( .A(n3728), .A(n3728_n), .B(n3796), .B(n3796_n), .Y(n3349_n), .Y(n3349) );
 NAND2X1TS U2760 ( .A(n3799), .A(n3799_n), .B(n3800), .B(n3800_n), .Y(n3798_n), .Y(n3798) );
 NAND2X1TS U2761 ( .A(n3062), .A(n3062_n), .B(n3801), .B(n3801_n), .Y(n3800_n), .Y(n3800) );
 NAND2X1TS U2762 ( .A(n3706), .A(n3706_n), .B(n3086), .B(n3086_n), .Y(n3801_n), .Y(n3801) );
 NAND2X1TS U2763 ( .A(n3008), .A(n3008_n), .B(n3257), .B(n3257_n), .Y(n3799_n), .Y(n3799) );
 NAND2X1TS U2764 ( .A(n3805), .A(n3805_n), .B(n3806), .B(n3806_n), .Y(n3793_n), .Y(n3793) );
 NAND2X1TS U2765 ( .A(n3121), .A(n3121_n), .B(n3028), .B(n3028_n), .Y(n3758_n), .Y(n3758) );
 NAND2X1TS U2766 ( .A(n3811), .A(n3811_n), .B(n3312), .B(n3312_n), .Y(n3810_n), .Y(n3810) );
 NAND2X1TS U2767 ( .A(n3025), .A(n3025_n), .B(n3457), .B(n3457_n), .Y(n3312_n), .Y(n3312) );
 NAND2X1TS U2768 ( .A(n3863), .A(n3863_n), .B(n3784), .B(n3784_n), .Y(n3175_n), .Y(n3175) );
 NAND2X1TS U2769 ( .A(n3043), .A(n3043_n), .B(n3298), .B(n3298_n), .Y(n3811_n), .Y(n3811) );
 NAND2X1TS U2770 ( .A(n3813), .A(n3813_n), .B(n3595), .B(n3595_n), .Y(n3809_n), .Y(n3809) );
 NAND2X1TS U2771 ( .A(n3083), .A(n3083_n), .B(n2997), .B(n2997_n), .Y(n3595_n), .Y(n3595) );
 NAND2X1TS U2772 ( .A(n3115), .A(n3115_n), .B(n2966), .B(n2966_n), .Y(n3626_n), .Y(n3626) );
 NAND2X1TS U2773 ( .A(n3204), .A(n3204_n), .B(n3677), .B(n3677_n), .Y(n3127_n), .Y(n3127) );
 NAND2X1TS U2774 ( .A(n3680), .A(n3680_n), .B(n3391), .B(n3391_n), .Y(n3679_n), .Y(n3679) );
 NAND2X1TS U2775 ( .A(n3184), .A(n3184_n), .B(n3199), .B(n3199_n), .Y(n3391_n), .Y(n3391) );
 NAND2X1TS U2776 ( .A(n3117), .A(n3117_n), .B(n3148), .B(n3148_n), .Y(n3829_n), .Y(n3829) );
 NAND2X1TS U2777 ( .A(n3334), .A(n3334_n), .B(n3296), .B(n3296_n), .Y(n3682_n), .Y(n3682) );
 NAND2X1TS U2778 ( .A(n3071), .A(n3071_n), .B(n3066), .B(n3066_n), .Y(n3296_n), .Y(n3296) );
 NAND2X1TS U2779 ( .A(n3032), .A(n3032_n), .B(n3040), .B(n3040_n), .Y(n3334_n), .Y(n3334) );
 NAND2X1TS U2780 ( .A(n3313), .A(n3313_n), .B(n3683), .B(n3683_n), .Y(n3681_n), .Y(n3681) );
 NAND2X1TS U2781 ( .A(n3465), .A(n3465_n), .B(n3062), .B(n3062_n), .Y(n3683_n), .Y(n3683) );
 NAND2X1TS U2782 ( .A(n3110), .A(n3110_n), .B(n3859), .B(n3859_n), .Y(n3510_n), .Y(n3510) );
 NAND2X1TS U2783 ( .A(n2998), .A(n2998_n), .B(n3044), .B(n3044_n), .Y(n3313_n), .Y(n3313) );
 NAND2X1TS U2784 ( .A(n3684), .A(n3684_n), .B(n3685), .B(n3685_n), .Y(n3678_n), .Y(n3678) );
 NAND2X1TS U2785 ( .A(n3028), .A(n3028_n), .B(n3686), .B(n3686_n), .Y(n3685_n), .Y(n3685) );
 NAND2X1TS U2786 ( .A(n3575), .A(n3575_n), .B(n3005), .B(n3005_n), .Y(n3686_n), .Y(n3686) );
 NAND2X1TS U2787 ( .A(n3689), .A(n3689_n), .B(n3690), .B(n3690_n), .Y(n3688_n), .Y(n3688) );
 NAND2X1TS U2788 ( .A(n3007), .A(n3007_n), .B(n3396), .B(n3396_n), .Y(n3690_n), .Y(n3690) );
 NAND2X1TS U2789 ( .A(n3156), .A(n3156_n), .B(n3443), .B(n3443_n), .Y(n3396_n), .Y(n3396) );
 NAND2X1TS U2790 ( .A(n2971), .A(n2971_n), .B(n3789), .B(n3789_n), .Y(n3692_n), .Y(n3692) );
 NAND2X1TS U2791 ( .A(n3693), .A(n3693_n), .B(n3694), .B(n3694_n), .Y(n3687_n), .Y(n3687) );
 NAND2X1TS U2792 ( .A(n3065), .A(n3065_n), .B(n3449), .B(n3449_n), .Y(n3694_n), .Y(n3694) );
 NAND2X1TS U2793 ( .A(n3699), .A(n3699_n), .B(n3700), .B(n3700_n), .Y(n3698_n), .Y(n3698) );
 NAND2X1TS U2794 ( .A(n3022), .A(n3022_n), .B(n3701), .B(n3701_n), .Y(n3700_n), .Y(n3700) );
 NAND2X1TS U2795 ( .A(n3551), .A(n3551_n), .B(n2987), .B(n2987_n), .Y(n3701_n), .Y(n3701) );
 NAND2X1TS U2796 ( .A(n3443), .A(n3443_n), .B(n3535), .B(n3535_n), .Y(n3147_n), .Y(n3147) );
 NAND2X1TS U2797 ( .A(n3122), .A(n3122_n), .B(n2996), .B(n2996_n), .Y(n3535_n), .Y(n3535) );
 NAND2X1TS U2798 ( .A(n3704), .A(n3704_n), .B(n3381), .B(n3381_n), .Y(n3703_n), .Y(n3703) );
 NAND2X1TS U2799 ( .A(n3417), .A(n3417_n), .B(n3198), .B(n3198_n), .Y(n3381_n), .Y(n3381) );
 NAND2X1TS U2800 ( .A(n3718), .A(n3718_n), .B(n3785), .B(n3785_n), .Y(n3291_n), .Y(n3291) );
 NAND2X1TS U2801 ( .A(n3105), .A(n3105_n), .B(n3106), .B(n3106_n), .Y(n3869_n), .Y(n3869) );
 NAND2X1TS U2802 ( .A(n3784), .A(n3784_n), .B(n3785), .B(n3785_n), .Y(n3319_n), .Y(n3319) );
 NAND2X1TS U2803 ( .A(n3115), .A(n3115_n), .B(n2964), .B(n2964_n), .Y(n3540_n), .Y(n3540) );
 NAND2X1TS U2804 ( .A(n3707), .A(n3707_n), .B(n3708), .B(n3708_n), .Y(n3697_n), .Y(n3697) );
 NAND2X1TS U2805 ( .A(n3711), .A(n3711_n), .B(n3712), .B(n3712_n), .Y(n3710_n), .Y(n3710) );
 NAND2X1TS U2806 ( .A(n3077), .A(n3077_n), .B(n3140), .B(n3140_n), .Y(n3712_n), .Y(n3712) );
 NAND2X1TS U2807 ( .A(n2978), .A(n2978_n), .B(n2985), .B(n2985_n), .Y(n3443_n), .Y(n3443) );
 NAND2X1TS U2808 ( .A(n2966), .A(n2966_n), .B(n3030), .B(n3030_n), .Y(n3235_n), .Y(n3235) );
 NAND2X1TS U2809 ( .A(n3859), .A(n3859_n), .B(n3109), .B(n3109_n), .Y(n3265_n), .Y(n3265) );
 NAND2X1TS U2810 ( .A(n2958), .A(n2958_n), .B(n3141), .B(n3141_n), .Y(n3711_n), .Y(n3711) );
 NAND2X1TS U2811 ( .A(n3055), .A(n3055_n), .B(n3316), .B(n3316_n), .Y(n3141_n), .Y(n3141) );
 NAND2X1TS U2812 ( .A(n2980), .A(n2980_n), .B(n3029), .B(n3029_n), .Y(n3764_n), .Y(n3764) );
 NAND2X1TS U2813 ( .A(n3189), .A(n3189_n), .B(n3715), .B(n3715_n), .Y(n3714_n), .Y(n3714) );
 NAND2X1TS U2814 ( .A(n3654), .A(n3654_n), .B(n3716), .B(n3716_n), .Y(n3715_n), .Y(n3715) );
 NAND2X1TS U2815 ( .A(n3713), .A(n3713_n), .B(n3717), .B(n3717_n), .Y(n3716_n), .Y(n3716) );
 NAND2X1TS U2816 ( .A(n3119), .A(n3119_n), .B(n3718), .B(n3718_n), .Y(n3717_n), .Y(n3717) );
 NAND2X1TS U2817 ( .A(n2977), .A(n2977_n), .B(n2971), .B(n2971_n), .Y(n3858_n), .Y(n3858) );
 NAND2X1TS U2818 ( .A(n3114), .A(n3114_n), .B(n2995), .B(n2995_n), .Y(n3549_n), .Y(n3549) );
 NAND2X1TS U2819 ( .A(n3082), .A(n3082_n), .B(n3608), .B(n3608_n), .Y(n3189_n), .Y(n3189) );
 NAND2X1TS U2820 ( .A(n3123), .A(n3123_n), .B(n3000), .B(n3000_n), .Y(n3720_n), .Y(n3720) );
 NAND2X1TS U2821 ( .A(n3113), .A(n3113_n), .B(n3027), .B(n3027_n), .Y(n3550_n), .Y(n3550) );
 NAND2X1TS U2822 ( .A(n3110), .A(n3110_n), .B(n3876), .B(n3876_n), .Y(n3173_n), .Y(n3173) );
endmodule

