`timescale 1ns/100ps

module beta_alu_tb;

reg clock = 0;
integer dut_error = 0;

reg  [31:0] a;
reg  [31:0] b;
reg   [5:0] fn;
wire [31:0] y;

// -------------------------------------------------------
// CLOCK GENERATION
// -------------------------------------------------------

always begin
	clock=0; #4;  // 125 MHz
	clock=1; #4;
end

// -------------------------------------------------------
// INITIALIZATION
// -------------------------------------------------------

initial begin
	if ($test$plusargs("vcd")) begin
		$dumpfile ("beta_alu_tb.vcd");
		$dumpvars (5, beta_alu_tb, dut);
	end
end

// -------------------------------------------------------
// TEST CASES
// -------------------------------------------------------

task test_case;
    input [69:0] inputs;
    input [34:0] expected_output;
	input integer line;
    begin
        {fn, a, b} <= inputs;
        @(posedge clock)
        if ({y, dut.z, dut.v, dut.n} == expected_output) begin
            $display("pass:  fn=%02x, a=%08x, b=%08x => y=%08x, zvn=%01x",
                     inputs[69:64], inputs[63:32], inputs[31:0],
                     y, {dut.z, dut.v, dut.n});
        end else begin
            $display("FAIL:  fn=%02x, a=%08x, b=%02x => y=%08x, zvn=%01x (expected %08x, %01x)",
                     inputs[69:64], inputs[63:32], inputs[31:0],
                     y, {dut.z, dut.v, dut.n},
                     expected_output[34:3], expected_output[2:0]);
			$error("");
			$display("       test_case at line %d", line);
			dut_error = dut_error + 1;
        end
    end
endtask

initial begin
	@(posedge clock);
	$display("");
	test_case({6'b100010, 32'b11111111000000001111111100000000, 32'b11111111111111110000000000000000}, {32'b00000000000000001111111100000000, 3'b001}, `__LINE__); //   3: fn=F0010, a=0xff00ff00, b=0xffff0000, y=0x0000ff00
	test_case({6'b100001, 32'b11111111000000001111111100000000, 32'b11111111111111110000000000000000}, {32'b00000000000000000000000011111111, 3'b001}, `__LINE__); //   2: fn=F0001, a=0xff00ff00, b=0xffff0000, y=0x000000ff
	test_case({6'b100011, 32'b11111111000000001111111100000000, 32'b11111111111111110000000000000000}, {32'b00000000000000001111111111111111, 3'b001}, `__LINE__); //   4: fn=F0011, a=0xff00ff00, b=0xffff0000, y=0x0000ffff
	test_case({6'b100100, 32'b11111111000000001111111100000000, 32'b11111111111111110000000000000000}, {32'b00000000111111110000000000000000, 3'b001}, `__LINE__); //   5: fn=F0100, a=0xff00ff00, b=0xffff0000, y=0x00ff0000
	test_case({6'b100101, 32'b11111111000000001111111100000000, 32'b11111111111111110000000000000000}, {32'b00000000111111110000000011111111, 3'b001}, `__LINE__); //   6: fn=F0101, a=0xff00ff00, b=0xffff0000, y=0x00ff00ff
	test_case({6'b100110, 32'b11111111000000001111111100000000, 32'b11111111111111110000000000000000}, {32'b00000000111111111111111100000000, 3'b001}, `__LINE__); //   7: fn=  XOR, a=0xff00ff00, b=0xffff0000, y=0x00ffff00
	test_case({6'b101000, 32'b11111111000000001111111100000000, 32'b11111111111111110000000000000000}, {32'b11111111000000000000000000000000, 3'b001}, `__LINE__); //   9: fn=  AND, a=0xff00ff00, b=0xffff0000, y=0xff000000
	test_case({6'b100111, 32'b11111111000000001111111100000000, 32'b11111111111111110000000000000000}, {32'b00000000111111111111111111111111, 3'b001}, `__LINE__); //   8: fn=F0111, a=0xff00ff00, b=0xffff0000, y=0x00ffffff
	test_case({6'b100000, 32'b11111111000000001111111100000000, 32'b11111111111111110000000000000000}, {32'b00000000000000000000000000000000, 3'b001}, `__LINE__); //   1: fn=F0000, a=0xff00ff00, b=0xffff0000, y=0x00000000
	test_case({6'b101001, 32'b11111111000000001111111100000000, 32'b11111111111111110000000000000000}, {32'b11111111000000000000000011111111, 3'b001}, `__LINE__); //  10: fn= XNOR, a=0xff00ff00, b=0xffff0000, y=0xff0000ff
	test_case({6'b101010, 32'b11111111000000001111111100000000, 32'b11111111111111110000000000000000}, {32'b11111111000000001111111100000000, 3'b001}, `__LINE__); //  11: fn=    A, a=0xff00ff00, b=0xffff0000, y=0xff00ff00
	test_case({6'b101011, 32'b11111111000000001111111100000000, 32'b11111111111111110000000000000000}, {32'b11111111000000001111111111111111, 3'b001}, `__LINE__); //  12: fn=F1011, a=0xff00ff00, b=0xffff0000, y=0xff00ffff
	test_case({6'b101100, 32'b11111111000000001111111100000000, 32'b11111111111111110000000000000000}, {32'b11111111111111110000000000000000, 3'b001}, `__LINE__); //  13: fn=F1100, a=0xff00ff00, b=0xffff0000, y=0xffff0000
	test_case({6'b101101, 32'b11111111000000001111111100000000, 32'b11111111111111110000000000000000}, {32'b11111111111111110000000011111111, 3'b001}, `__LINE__); //  14: fn=F1101, a=0xff00ff00, b=0xffff0000, y=0xffff00ff
	test_case({6'b101110, 32'b11111111000000001111111100000000, 32'b11111111111111110000000000000000}, {32'b11111111111111111111111100000000, 3'b001}, `__LINE__); //  15: fn=   OR, a=0xff00ff00, b=0xffff0000, y=0xffffff00
	test_case({6'b101111, 32'b11111111000000001111111100000000, 32'b11111111111111110000000000000000}, {32'b11111111111111111111111111111111, 3'b001}, `__LINE__); //  16: fn=F1111, a=0xff00ff00, b=0xffff0000, y=0xffffffff
	test_case({6'b110000, 32'b00000000000000000000000000000000, 32'b00000000000000000000000000000000}, {32'b00000000000000000000000000000000, 3'b100}, `__LINE__); //  17: fn=  SHL, a=0x00000000, b=0x00000000, y=0x00000000
	test_case({6'b110001, 32'b00000000000000000000000000000000, 32'b00000000000000000000000000000000}, {32'b00000000000000000000000000000000, 3'b100}, `__LINE__); //  18: fn=  SHR, a=0x00000000, b=0x00000000, y=0x00000000
	test_case({6'b110011, 32'b00000000000000000000000000000000, 32'b00000000000000000000000000000000}, {32'b00000000000000000000000000000000, 3'b100}, `__LINE__); //  19: fn=  SRA, a=0x00000000, b=0x00000000, y=0x00000000
	test_case({6'b110000, 32'b00000000000000000000000000000000, 32'b00000000000000000000000000000001}, {32'b00000000000000000000000000000000, 3'b000}, `__LINE__); //  20: fn=  SHL, a=0x00000000, b=0x00000001, y=0x00000000
	test_case({6'b110001, 32'b00000000000000000000000000000000, 32'b00000000000000000000000000000001}, {32'b00000000000000000000000000000000, 3'b001}, `__LINE__); //  21: fn=  SHR, a=0x00000000, b=0x00000001, y=0x00000000
	test_case({6'b110011, 32'b00000000000000000000000000000000, 32'b00000000000000000000000000000001}, {32'b00000000000000000000000000000000, 3'b001}, `__LINE__); //  22: fn=  SRA, a=0x00000000, b=0x00000001, y=0x00000000
	test_case({6'b110000, 32'b00000000000000000000000000000000, 32'b00000000000000000000000000000010}, {32'b00000000000000000000000000000000, 3'b000}, `__LINE__); //  23: fn=  SHL, a=0x00000000, b=0x00000002, y=0x00000000
	test_case({6'b110001, 32'b00000000000000000000000000000000, 32'b00000000000000000000000000000010}, {32'b00000000000000000000000000000000, 3'b001}, `__LINE__); //  24: fn=  SHR, a=0x00000000, b=0x00000002, y=0x00000000
	test_case({6'b110011, 32'b00000000000000000000000000000000, 32'b00000000000000000000000000000010}, {32'b00000000000000000000000000000000, 3'b001}, `__LINE__); //  25: fn=  SRA, a=0x00000000, b=0x00000002, y=0x00000000
	test_case({6'b110000, 32'b00000000000000000000000000000000, 32'b00000000000000000000000000000100}, {32'b00000000000000000000000000000000, 3'b000}, `__LINE__); //  26: fn=  SHL, a=0x00000000, b=0x00000004, y=0x00000000
	test_case({6'b110001, 32'b00000000000000000000000000000000, 32'b00000000000000000000000000000100}, {32'b00000000000000000000000000000000, 3'b001}, `__LINE__); //  27: fn=  SHR, a=0x00000000, b=0x00000004, y=0x00000000
	test_case({6'b110011, 32'b00000000000000000000000000000000, 32'b00000000000000000000000000000100}, {32'b00000000000000000000000000000000, 3'b001}, `__LINE__); //  28: fn=  SRA, a=0x00000000, b=0x00000004, y=0x00000000
	test_case({6'b110000, 32'b00000000000000000000000000000000, 32'b00000000000000000000000000001000}, {32'b00000000000000000000000000000000, 3'b000}, `__LINE__); //  29: fn=  SHL, a=0x00000000, b=0x00000008, y=0x00000000
	test_case({6'b110001, 32'b00000000000000000000000000000000, 32'b00000000000000000000000000001000}, {32'b00000000000000000000000000000000, 3'b001}, `__LINE__); //  30: fn=  SHR, a=0x00000000, b=0x00000008, y=0x00000000
	test_case({6'b110011, 32'b00000000000000000000000000000000, 32'b00000000000000000000000000001000}, {32'b00000000000000000000000000000000, 3'b001}, `__LINE__); //  31: fn=  SRA, a=0x00000000, b=0x00000008, y=0x00000000
	test_case({6'b110000, 32'b00000000000000000000000000000000, 32'b00000000000000000000000000010000}, {32'b00000000000000000000000000000000, 3'b000}, `__LINE__); //  32: fn=  SHL, a=0x00000000, b=0x00000010, y=0x00000000
	test_case({6'b110001, 32'b00000000000000000000000000000000, 32'b00000000000000000000000000010000}, {32'b00000000000000000000000000000000, 3'b001}, `__LINE__); //  33: fn=  SHR, a=0x00000000, b=0x00000010, y=0x00000000
	test_case({6'b110011, 32'b00000000000000000000000000000000, 32'b00000000000000000000000000010000}, {32'b00000000000000000000000000000000, 3'b001}, `__LINE__); //  34: fn=  SRA, a=0x00000000, b=0x00000010, y=0x00000000
	test_case({6'b110000, 32'b00000000000000000000000000000000, 32'b00000000000000000000000000011111}, {32'b00000000000000000000000000000000, 3'b000}, `__LINE__); //  35: fn=  SHL, a=0x00000000, b=0x0000001f, y=0x00000000
	test_case({6'b110001, 32'b00000000000000000000000000000000, 32'b00000000000000000000000000011111}, {32'b00000000000000000000000000000000, 3'b001}, `__LINE__); //  36: fn=  SHR, a=0x00000000, b=0x0000001f, y=0x00000000
	test_case({6'b110011, 32'b00000000000000000000000000000000, 32'b00000000000000000000000000011111}, {32'b00000000000000000000000000000000, 3'b001}, `__LINE__); //  37: fn=  SRA, a=0x00000000, b=0x0000001f, y=0x00000000
	test_case({6'b110000, 32'b00000000000000000000000000000001, 32'b00000000000000000000000000000000}, {32'b00000000000000000000000000000001, 3'b000}, `__LINE__); //  38: fn=  SHL, a=0x00000001, b=0x00000000, y=0x00000001
	test_case({6'b110001, 32'b00000000000000000000000000000001, 32'b00000000000000000000000000000000}, {32'b00000000000000000000000000000001, 3'b000}, `__LINE__); //  39: fn=  SHR, a=0x00000001, b=0x00000000, y=0x00000001
	test_case({6'b110011, 32'b00000000000000000000000000000001, 32'b00000000000000000000000000000000}, {32'b00000000000000000000000000000001, 3'b000}, `__LINE__); //  40: fn=  SRA, a=0x00000001, b=0x00000000, y=0x00000001
	test_case({6'b110000, 32'b00000000000000000000000000000001, 32'b00000000000000000000000000000001}, {32'b00000000000000000000000000000010, 3'b000}, `__LINE__); //  41: fn=  SHL, a=0x00000001, b=0x00000001, y=0x00000002
	test_case({6'b110001, 32'b00000000000000000000000000000001, 32'b00000000000000000000000000000001}, {32'b00000000000000000000000000000000, 3'b100}, `__LINE__); //  42: fn=  SHR, a=0x00000001, b=0x00000001, y=0x00000000
	test_case({6'b110011, 32'b00000000000000000000000000000001, 32'b00000000000000000000000000000001}, {32'b00000000000000000000000000000000, 3'b100}, `__LINE__); //  43: fn=  SRA, a=0x00000001, b=0x00000001, y=0x00000000
	test_case({6'b110000, 32'b00000000000000000000000000000001, 32'b00000000000000000000000000000010}, {32'b00000000000000000000000000000100, 3'b000}, `__LINE__); //  44: fn=  SHL, a=0x00000001, b=0x00000002, y=0x00000004
	test_case({6'b110001, 32'b00000000000000000000000000000001, 32'b00000000000000000000000000000010}, {32'b00000000000000000000000000000000, 3'b001}, `__LINE__); //  45: fn=  SHR, a=0x00000001, b=0x00000002, y=0x00000000
	test_case({6'b110011, 32'b00000000000000000000000000000001, 32'b00000000000000000000000000000010}, {32'b00000000000000000000000000000000, 3'b001}, `__LINE__); //  46: fn=  SRA, a=0x00000001, b=0x00000002, y=0x00000000
	test_case({6'b110000, 32'b00000000000000000000000000000001, 32'b00000000000000000000000000000100}, {32'b00000000000000000000000000010000, 3'b000}, `__LINE__); //  47: fn=  SHL, a=0x00000001, b=0x00000004, y=0x00000010
	test_case({6'b110001, 32'b00000000000000000000000000000001, 32'b00000000000000000000000000000100}, {32'b00000000000000000000000000000000, 3'b001}, `__LINE__); //  48: fn=  SHR, a=0x00000001, b=0x00000004, y=0x00000000
	test_case({6'b110011, 32'b00000000000000000000000000000001, 32'b00000000000000000000000000000100}, {32'b00000000000000000000000000000000, 3'b001}, `__LINE__); //  49: fn=  SRA, a=0x00000001, b=0x00000004, y=0x00000000
	test_case({6'b110000, 32'b00000000000000000000000000000001, 32'b00000000000000000000000000001000}, {32'b00000000000000000000000100000000, 3'b000}, `__LINE__); //  50: fn=  SHL, a=0x00000001, b=0x00000008, y=0x00000100
	test_case({6'b110001, 32'b00000000000000000000000000000001, 32'b00000000000000000000000000001000}, {32'b00000000000000000000000000000000, 3'b001}, `__LINE__); //  51: fn=  SHR, a=0x00000001, b=0x00000008, y=0x00000000
	test_case({6'b110011, 32'b00000000000000000000000000000001, 32'b00000000000000000000000000001000}, {32'b00000000000000000000000000000000, 3'b001}, `__LINE__); //  52: fn=  SRA, a=0x00000001, b=0x00000008, y=0x00000000
	test_case({6'b110000, 32'b00000000000000000000000000000001, 32'b00000000000000000000000000010000}, {32'b00000000000000010000000000000000, 3'b000}, `__LINE__); //  53: fn=  SHL, a=0x00000001, b=0x00000010, y=0x00010000
	test_case({6'b110001, 32'b00000000000000000000000000000001, 32'b00000000000000000000000000010000}, {32'b00000000000000000000000000000000, 3'b001}, `__LINE__); //  54: fn=  SHR, a=0x00000001, b=0x00000010, y=0x00000000
	test_case({6'b110011, 32'b00000000000000000000000000000001, 32'b00000000000000000000000000010000}, {32'b00000000000000000000000000000000, 3'b001}, `__LINE__); //  55: fn=  SRA, a=0x00000001, b=0x00000010, y=0x00000000
	test_case({6'b110000, 32'b00000000000000000000000000000001, 32'b00000000000000000000000000011111}, {32'b10000000000000000000000000000000, 3'b000}, `__LINE__); //  56: fn=  SHL, a=0x00000001, b=0x0000001f, y=0x80000000
	test_case({6'b110001, 32'b00000000000000000000000000000001, 32'b00000000000000000000000000011111}, {32'b00000000000000000000000000000000, 3'b001}, `__LINE__); //  57: fn=  SHR, a=0x00000001, b=0x0000001f, y=0x00000000
	test_case({6'b110011, 32'b00000000000000000000000000000001, 32'b00000000000000000000000000011111}, {32'b00000000000000000000000000000000, 3'b001}, `__LINE__); //  58: fn=  SRA, a=0x00000001, b=0x0000001f, y=0x00000000
	test_case({6'b110000, 32'b11111111111111111111111111111111, 32'b00000000000000000000000000000000}, {32'b11111111111111111111111111111111, 3'b001}, `__LINE__); //  59: fn=  SHL, a=0xffffffff, b=0x00000000, y=0xffffffff
	test_case({6'b110001, 32'b11111111111111111111111111111111, 32'b00000000000000000000000000000000}, {32'b11111111111111111111111111111111, 3'b001}, `__LINE__); //  60: fn=  SHR, a=0xffffffff, b=0x00000000, y=0xffffffff
	test_case({6'b110011, 32'b11111111111111111111111111111111, 32'b00000000000000000000000000000000}, {32'b11111111111111111111111111111111, 3'b001}, `__LINE__); //  61: fn=  SRA, a=0xffffffff, b=0x00000000, y=0xffffffff
	test_case({6'b110000, 32'b11111111111111111111111111111111, 32'b00000000000000000000000000000001}, {32'b11111111111111111111111111111110, 3'b100}, `__LINE__); //  62: fn=  SHL, a=0xffffffff, b=0x00000001, y=0xfffffffe
	test_case({6'b110001, 32'b11111111111111111111111111111111, 32'b00000000000000000000000000000001}, {32'b01111111111111111111111111111111, 3'b001}, `__LINE__); //  63: fn=  SHR, a=0xffffffff, b=0x00000001, y=0x7fffffff
	test_case({6'b110011, 32'b11111111111111111111111111111111, 32'b00000000000000000000000000000001}, {32'b11111111111111111111111111111111, 3'b001}, `__LINE__); //  64: fn=  SRA, a=0xffffffff, b=0x00000001, y=0xffffffff
	test_case({6'b110000, 32'b11111111111111111111111111111111, 32'b00000000000000000000000000000010}, {32'b11111111111111111111111111111100, 3'b000}, `__LINE__); //  65: fn=  SHL, a=0xffffffff, b=0x00000002, y=0xfffffffc
	test_case({6'b110001, 32'b11111111111111111111111111111111, 32'b00000000000000000000000000000010}, {32'b00111111111111111111111111111111, 3'b001}, `__LINE__); //  66: fn=  SHR, a=0xffffffff, b=0x00000002, y=0x3fffffff
	test_case({6'b110011, 32'b11111111111111111111111111111111, 32'b00000000000000000000000000000010}, {32'b11111111111111111111111111111111, 3'b001}, `__LINE__); //  67: fn=  SRA, a=0xffffffff, b=0x00000002, y=0xffffffff
	test_case({6'b110000, 32'b11111111111111111111111111111111, 32'b00000000000000000000000000000100}, {32'b11111111111111111111111111110000, 3'b000}, `__LINE__); //  68: fn=  SHL, a=0xffffffff, b=0x00000004, y=0xfffffff0
	test_case({6'b110001, 32'b11111111111111111111111111111111, 32'b00000000000000000000000000000100}, {32'b00001111111111111111111111111111, 3'b001}, `__LINE__); //  69: fn=  SHR, a=0xffffffff, b=0x00000004, y=0x0fffffff
	test_case({6'b110011, 32'b11111111111111111111111111111111, 32'b00000000000000000000000000000100}, {32'b11111111111111111111111111111111, 3'b001}, `__LINE__); //  70: fn=  SRA, a=0xffffffff, b=0x00000004, y=0xffffffff
	test_case({6'b110000, 32'b11111111111111111111111111111111, 32'b00000000000000000000000000001000}, {32'b11111111111111111111111100000000, 3'b000}, `__LINE__); //  71: fn=  SHL, a=0xffffffff, b=0x00000008, y=0xffffff00
	test_case({6'b110001, 32'b11111111111111111111111111111111, 32'b00000000000000000000000000001000}, {32'b00000000111111111111111111111111, 3'b001}, `__LINE__); //  72: fn=  SHR, a=0xffffffff, b=0x00000008, y=0x00ffffff
	test_case({6'b110011, 32'b11111111111111111111111111111111, 32'b00000000000000000000000000001000}, {32'b11111111111111111111111111111111, 3'b001}, `__LINE__); //  73: fn=  SRA, a=0xffffffff, b=0x00000008, y=0xffffffff
	test_case({6'b110000, 32'b11111111111111111111111111111111, 32'b00000000000000000000000000010000}, {32'b11111111111111110000000000000000, 3'b000}, `__LINE__); //  74: fn=  SHL, a=0xffffffff, b=0x00000010, y=0xffff0000
	test_case({6'b110001, 32'b11111111111111111111111111111111, 32'b00000000000000000000000000010000}, {32'b00000000000000001111111111111111, 3'b001}, `__LINE__); //  75: fn=  SHR, a=0xffffffff, b=0x00000010, y=0x0000ffff
	test_case({6'b110011, 32'b11111111111111111111111111111111, 32'b00000000000000000000000000010000}, {32'b11111111111111111111111111111111, 3'b001}, `__LINE__); //  76: fn=  SRA, a=0xffffffff, b=0x00000010, y=0xffffffff
	test_case({6'b110000, 32'b11111111111111111111111111111111, 32'b00000000000000000000000000011111}, {32'b10000000000000000000000000000000, 3'b000}, `__LINE__); //  77: fn=  SHL, a=0xffffffff, b=0x0000001f, y=0x80000000
	test_case({6'b110001, 32'b11111111111111111111111111111111, 32'b00000000000000000000000000011111}, {32'b00000000000000000000000000000001, 3'b001}, `__LINE__); //  78: fn=  SHR, a=0xffffffff, b=0x0000001f, y=0x00000001
	test_case({6'b110011, 32'b11111111111111111111111111111111, 32'b00000000000000000000000000011111}, {32'b11111111111111111111111111111111, 3'b001}, `__LINE__); //  79: fn=  SRA, a=0xffffffff, b=0x0000001f, y=0xffffffff
	test_case({6'b110000, 32'b00010010001101000101011001111000, 32'b00000000000000000000000000000000}, {32'b00010010001101000101011001111000, 3'b000}, `__LINE__); //  80: fn=  SHL, a=0x12345678, b=0x00000000, y=0x12345678
	test_case({6'b110001, 32'b00010010001101000101011001111000, 32'b00000000000000000000000000000000}, {32'b00010010001101000101011001111000, 3'b000}, `__LINE__); //  81: fn=  SHR, a=0x12345678, b=0x00000000, y=0x12345678
	test_case({6'b110011, 32'b00010010001101000101011001111000, 32'b00000000000000000000000000000000}, {32'b00010010001101000101011001111000, 3'b000}, `__LINE__); //  82: fn=  SRA, a=0x12345678, b=0x00000000, y=0x12345678
	test_case({6'b110000, 32'b00010010001101000101011001111000, 32'b00000000000000000000000000000001}, {32'b00100100011010001010110011110000, 3'b000}, `__LINE__); //  83: fn=  SHL, a=0x12345678, b=0x00000001, y=0x2468acf0
	test_case({6'b110001, 32'b00010010001101000101011001111000, 32'b00000000000000000000000000000001}, {32'b00001001000110100010101100111100, 3'b000}, `__LINE__); //  84: fn=  SHR, a=0x12345678, b=0x00000001, y=0x091a2b3c
	test_case({6'b110011, 32'b00010010001101000101011001111000, 32'b00000000000000000000000000000001}, {32'b00001001000110100010101100111100, 3'b000}, `__LINE__); //  85: fn=  SRA, a=0x12345678, b=0x00000001, y=0x091a2b3c
	test_case({6'b110000, 32'b00010010001101000101011001111000, 32'b00000000000000000000000000000010}, {32'b01001000110100010101100111100000, 3'b000}, `__LINE__); //  86: fn=  SHL, a=0x12345678, b=0x00000002, y=0x48d159e0
	test_case({6'b110001, 32'b00010010001101000101011001111000, 32'b00000000000000000000000000000010}, {32'b00000100100011010001010110011110, 3'b000}, `__LINE__); //  87: fn=  SHR, a=0x12345678, b=0x00000002, y=0x048d159e
	test_case({6'b110011, 32'b00010010001101000101011001111000, 32'b00000000000000000000000000000010}, {32'b00000100100011010001010110011110, 3'b000}, `__LINE__); //  88: fn=  SRA, a=0x12345678, b=0x00000002, y=0x048d159e
	test_case({6'b110000, 32'b00010010001101000101011001111000, 32'b00000000000000000000000000000100}, {32'b00100011010001010110011110000000, 3'b000}, `__LINE__); //  89: fn=  SHL, a=0x12345678, b=0x00000004, y=0x23456780
	test_case({6'b110001, 32'b00010010001101000101011001111000, 32'b00000000000000000000000000000100}, {32'b00000001001000110100010101100111, 3'b000}, `__LINE__); //  90: fn=  SHR, a=0x12345678, b=0x00000004, y=0x01234567
	test_case({6'b110011, 32'b00010010001101000101011001111000, 32'b00000000000000000000000000000100}, {32'b00000001001000110100010101100111, 3'b000}, `__LINE__); //  91: fn=  SRA, a=0x12345678, b=0x00000004, y=0x01234567
	test_case({6'b110000, 32'b00010010001101000101011001111000, 32'b00000000000000000000000000001000}, {32'b00110100010101100111100000000000, 3'b000}, `__LINE__); //  92: fn=  SHL, a=0x12345678, b=0x00000008, y=0x34567800
	test_case({6'b110001, 32'b00010010001101000101011001111000, 32'b00000000000000000000000000001000}, {32'b00000000000100100011010001010110, 3'b000}, `__LINE__); //  93: fn=  SHR, a=0x12345678, b=0x00000008, y=0x00123456
	test_case({6'b110011, 32'b00010010001101000101011001111000, 32'b00000000000000000000000000001000}, {32'b00000000000100100011010001010110, 3'b000}, `__LINE__); //  94: fn=  SRA, a=0x12345678, b=0x00000008, y=0x00123456
	test_case({6'b110000, 32'b00010010001101000101011001111000, 32'b00000000000000000000000000010000}, {32'b01010110011110000000000000000000, 3'b000}, `__LINE__); //  95: fn=  SHL, a=0x12345678, b=0x00000010, y=0x56780000
	test_case({6'b110001, 32'b00010010001101000101011001111000, 32'b00000000000000000000000000010000}, {32'b00000000000000000001001000110100, 3'b000}, `__LINE__); //  96: fn=  SHR, a=0x12345678, b=0x00000010, y=0x00001234
	test_case({6'b110011, 32'b00010010001101000101011001111000, 32'b00000000000000000000000000010000}, {32'b00000000000000000001001000110100, 3'b000}, `__LINE__); //  97: fn=  SRA, a=0x12345678, b=0x00000010, y=0x00001234
	test_case({6'b110000, 32'b00010010001101000101011001111000, 32'b00000000000000000000000000011111}, {32'b00000000000000000000000000000000, 3'b000}, `__LINE__); //  98: fn=  SHL, a=0x12345678, b=0x0000001f, y=0x00000000
	test_case({6'b110001, 32'b00010010001101000101011001111000, 32'b00000000000000000000000000011111}, {32'b00000000000000000000000000000000, 3'b000}, `__LINE__); //  99: fn=  SHR, a=0x12345678, b=0x0000001f, y=0x00000000
	test_case({6'b110011, 32'b00010010001101000101011001111000, 32'b00000000000000000000000000011111}, {32'b00000000000000000000000000000000, 3'b000}, `__LINE__); // 100: fn=  SRA, a=0x12345678, b=0x0000001f, y=0x00000000
	test_case({6'b110000, 32'b11111110110111001010101110011000, 32'b00000000000000000000000000000000}, {32'b11111110110111001010101110011000, 3'b001}, `__LINE__); // 101: fn=  SHL, a=0xfedcab98, b=0x00000000, y=0xfedcab98
	test_case({6'b110001, 32'b11111110110111001010101110011000, 32'b00000000000000000000000000000000}, {32'b11111110110111001010101110011000, 3'b001}, `__LINE__); // 102: fn=  SHR, a=0xfedcab98, b=0x00000000, y=0xfedcab98
	test_case({6'b110011, 32'b11111110110111001010101110011000, 32'b00000000000000000000000000000000}, {32'b11111110110111001010101110011000, 3'b001}, `__LINE__); // 103: fn=  SRA, a=0xfedcab98, b=0x00000000, y=0xfedcab98
	test_case({6'b110000, 32'b11111110110111001010101110011000, 32'b00000000000000000000000000000001}, {32'b11111101101110010101011100110000, 3'b001}, `__LINE__); // 104: fn=  SHL, a=0xfedcab98, b=0x00000001, y=0xfdb95730
	test_case({6'b110001, 32'b11111110110111001010101110011000, 32'b00000000000000000000000000000001}, {32'b01111111011011100101010111001100, 3'b001}, `__LINE__); // 105: fn=  SHR, a=0xfedcab98, b=0x00000001, y=0x7f6e55cc
	test_case({6'b110011, 32'b11111110110111001010101110011000, 32'b00000000000000000000000000000001}, {32'b11111111011011100101010111001100, 3'b001}, `__LINE__); // 106: fn=  SRA, a=0xfedcab98, b=0x00000001, y=0xff6e55cc
	test_case({6'b110000, 32'b11111110110111001010101110011000, 32'b00000000000000000000000000000010}, {32'b11111011011100101010111001100000, 3'b001}, `__LINE__); // 107: fn=  SHL, a=0xfedcab98, b=0x00000002, y=0xfb72ae60
	test_case({6'b110001, 32'b11111110110111001010101110011000, 32'b00000000000000000000000000000010}, {32'b00111111101101110010101011100110, 3'b001}, `__LINE__); // 108: fn=  SHR, a=0xfedcab98, b=0x00000002, y=0x3fb72ae6
	test_case({6'b110011, 32'b11111110110111001010101110011000, 32'b00000000000000000000000000000010}, {32'b11111111101101110010101011100110, 3'b001}, `__LINE__); // 109: fn=  SRA, a=0xfedcab98, b=0x00000002, y=0xffb72ae6
	test_case({6'b110000, 32'b11111110110111001010101110011000, 32'b00000000000000000000000000000100}, {32'b11101101110010101011100110000000, 3'b001}, `__LINE__); // 110: fn=  SHL, a=0xfedcab98, b=0x00000004, y=0xedcab980
	test_case({6'b110001, 32'b11111110110111001010101110011000, 32'b00000000000000000000000000000100}, {32'b00001111111011011100101010111001, 3'b001}, `__LINE__); // 111: fn=  SHR, a=0xfedcab98, b=0x00000004, y=0x0fedcab9
	test_case({6'b110011, 32'b11111110110111001010101110011000, 32'b00000000000000000000000000000100}, {32'b11111111111011011100101010111001, 3'b001}, `__LINE__); // 112: fn=  SRA, a=0xfedcab98, b=0x00000004, y=0xffedcab9
	test_case({6'b110000, 32'b11111110110111001010101110011000, 32'b00000000000000000000000000001000}, {32'b11011100101010111001100000000000, 3'b001}, `__LINE__); // 113: fn=  SHL, a=0xfedcab98, b=0x00000008, y=0xdcab9800
	test_case({6'b110001, 32'b11111110110111001010101110011000, 32'b00000000000000000000000000001000}, {32'b00000000111111101101110010101011, 3'b001}, `__LINE__); // 114: fn=  SHR, a=0xfedcab98, b=0x00000008, y=0x00fedcab
	test_case({6'b110011, 32'b11111110110111001010101110011000, 32'b00000000000000000000000000001000}, {32'b11111111111111101101110010101011, 3'b001}, `__LINE__); // 115: fn=  SRA, a=0xfedcab98, b=0x00000008, y=0xfffedcab
	test_case({6'b110000, 32'b11111110110111001010101110011000, 32'b00000000000000000000000000010000}, {32'b10101011100110000000000000000000, 3'b001}, `__LINE__); // 116: fn=  SHL, a=0xfedcab98, b=0x00000010, y=0xab980000
	test_case({6'b110001, 32'b11111110110111001010101110011000, 32'b00000000000000000000000000010000}, {32'b00000000000000001111111011011100, 3'b001}, `__LINE__); // 117: fn=  SHR, a=0xfedcab98, b=0x00000010, y=0x0000fedc
	test_case({6'b110011, 32'b11111110110111001010101110011000, 32'b00000000000000000000000000010000}, {32'b11111111111111111111111011011100, 3'b001}, `__LINE__); // 118: fn=  SRA, a=0xfedcab98, b=0x00000010, y=0xfffffedc
	test_case({6'b110000, 32'b11111110110111001010101110011000, 32'b00000000000000000000000000011111}, {32'b00000000000000000000000000000000, 3'b001}, `__LINE__); // 119: fn=  SHL, a=0xfedcab98, b=0x0000001f, y=0x00000000
	test_case({6'b110001, 32'b11111110110111001010101110011000, 32'b00000000000000000000000000011111}, {32'b00000000000000000000000000000001, 3'b001}, `__LINE__); // 120: fn=  SHR, a=0xfedcab98, b=0x0000001f, y=0x00000001
	test_case({6'b110011, 32'b11111110110111001010101110011000, 32'b00000000000000000000000000011111}, {32'b11111111111111111111111111111111, 3'b001}, `__LINE__); // 121: fn=  SRA, a=0xfedcab98, b=0x0000001f, y=0xffffffff
	test_case({6'b010000, 32'b00000000000000000000000000000000, 32'b00000000000000000000000000000000}, {32'b00000000000000000000000000000000, 3'b100}, `__LINE__); // 122: fn=  ADD, a=0x00000000, b=0x00000000, y=0x00000000
	test_case({6'b010000, 32'b00000000000000000000000000000000, 32'b00000000000000000000000000000001}, {32'b00000000000000000000000000000001, 3'b000}, `__LINE__); // 123: fn=  ADD, a=0x00000000, b=0x00000001, y=0x00000001
	test_case({6'b010000, 32'b00000000000000000000000000000000, 32'b11111111111111111111111111111111}, {32'b11111111111111111111111111111111, 3'b001}, `__LINE__); // 124: fn=  ADD, a=0x00000000, b=0x-0000001, y=0xffffffff
	test_case({6'b010000, 32'b00000000000000000000000000000000, 32'b10101010101010101010101010101010}, {32'b10101010101010101010101010101010, 3'b001}, `__LINE__); // 125: fn=  ADD, a=0x00000000, b=0xaaaaaaaa, y=0xaaaaaaaa
	test_case({6'b010000, 32'b00000000000000000000000000000000, 32'b01010101010101010101010101010101}, {32'b01010101010101010101010101010101, 3'b000}, `__LINE__); // 126: fn=  ADD, a=0x00000000, b=0x55555555, y=0x55555555
	test_case({6'b010000, 32'b00000000000000000000000000000001, 32'b00000000000000000000000000000000}, {32'b00000000000000000000000000000001, 3'b000}, `__LINE__); // 127: fn=  ADD, a=0x00000001, b=0x00000000, y=0x00000001
	test_case({6'b010000, 32'b00000000000000000000000000000001, 32'b00000000000000000000000000000001}, {32'b00000000000000000000000000000010, 3'b000}, `__LINE__); // 128: fn=  ADD, a=0x00000001, b=0x00000001, y=0x00000002
	test_case({6'b010000, 32'b00000000000000000000000000000001, 32'b11111111111111111111111111111111}, {32'b00000000000000000000000000000000, 3'b100}, `__LINE__); // 129: fn=  ADD, a=0x00000001, b=0x-0000001, y=0x00000000
	test_case({6'b010000, 32'b00000000000000000000000000000001, 32'b10101010101010101010101010101010}, {32'b10101010101010101010101010101011, 3'b001}, `__LINE__); // 130: fn=  ADD, a=0x00000001, b=0xaaaaaaaa, y=0xaaaaaaab
	test_case({6'b010000, 32'b00000000000000000000000000000001, 32'b01010101010101010101010101010101}, {32'b01010101010101010101010101010110, 3'b000}, `__LINE__); // 131: fn=  ADD, a=0x00000001, b=0x55555555, y=0x55555556
	test_case({6'b010000, 32'b11111111111111111111111111111111, 32'b00000000000000000000000000000000}, {32'b11111111111111111111111111111111, 3'b001}, `__LINE__); // 132: fn=  ADD, a=0x-0000001, b=0x00000000, y=0xffffffff
	test_case({6'b010000, 32'b11111111111111111111111111111111, 32'b00000000000000000000000000000001}, {32'b00000000000000000000000000000000, 3'b100}, `__LINE__); // 133: fn=  ADD, a=0x-0000001, b=0x00000001, y=0x00000000
	test_case({6'b010000, 32'b11111111111111111111111111111111, 32'b11111111111111111111111111111111}, {32'b11111111111111111111111111111110, 3'b001}, `__LINE__); // 134: fn=  ADD, a=0x-0000001, b=0x-0000001, y=0xfffffffe
	test_case({6'b010000, 32'b11111111111111111111111111111111, 32'b10101010101010101010101010101010}, {32'b10101010101010101010101010101001, 3'b001}, `__LINE__); // 135: fn=  ADD, a=0x-0000001, b=0xaaaaaaaa, y=0xaaaaaaa9
	test_case({6'b010000, 32'b11111111111111111111111111111111, 32'b01010101010101010101010101010101}, {32'b01010101010101010101010101010100, 3'b000}, `__LINE__); // 136: fn=  ADD, a=0x-0000001, b=0x55555555, y=0x55555554
	test_case({6'b010000, 32'b10101010101010101010101010101010, 32'b00000000000000000000000000000000}, {32'b10101010101010101010101010101010, 3'b001}, `__LINE__); // 137: fn=  ADD, a=0xaaaaaaaa, b=0x00000000, y=0xaaaaaaaa
	test_case({6'b010000, 32'b10101010101010101010101010101010, 32'b00000000000000000000000000000001}, {32'b10101010101010101010101010101011, 3'b001}, `__LINE__); // 138: fn=  ADD, a=0xaaaaaaaa, b=0x00000001, y=0xaaaaaaab
	test_case({6'b010000, 32'b10101010101010101010101010101010, 32'b11111111111111111111111111111111}, {32'b10101010101010101010101010101001, 3'b001}, `__LINE__); // 139: fn=  ADD, a=0xaaaaaaaa, b=0x-0000001, y=0xaaaaaaa9
	test_case({6'b010000, 32'b10101010101010101010101010101010, 32'b10101010101010101010101010101010}, {32'b01010101010101010101010101010100, 3'b010}, `__LINE__); // 140: fn=  ADD, a=0xaaaaaaaa, b=0xaaaaaaaa, y=0x55555554
	test_case({6'b010000, 32'b10101010101010101010101010101010, 32'b01010101010101010101010101010101}, {32'b11111111111111111111111111111111, 3'b001}, `__LINE__); // 141: fn=  ADD, a=0xaaaaaaaa, b=0x55555555, y=0xffffffff
	test_case({6'b010000, 32'b01010101010101010101010101010101, 32'b00000000000000000000000000000000}, {32'b01010101010101010101010101010101, 3'b000}, `__LINE__); // 142: fn=  ADD, a=0x55555555, b=0x00000000, y=0x55555555
	test_case({6'b010000, 32'b01010101010101010101010101010101, 32'b00000000000000000000000000000001}, {32'b01010101010101010101010101010110, 3'b000}, `__LINE__); // 143: fn=  ADD, a=0x55555555, b=0x00000001, y=0x55555556
	test_case({6'b010000, 32'b01010101010101010101010101010101, 32'b11111111111111111111111111111111}, {32'b01010101010101010101010101010100, 3'b000}, `__LINE__); // 144: fn=  ADD, a=0x55555555, b=0x-0000001, y=0x55555554
	test_case({6'b010000, 32'b01010101010101010101010101010101, 32'b10101010101010101010101010101010}, {32'b11111111111111111111111111111111, 3'b001}, `__LINE__); // 145: fn=  ADD, a=0x55555555, b=0xaaaaaaaa, y=0xffffffff
	test_case({6'b010000, 32'b01010101010101010101010101010101, 32'b01010101010101010101010101010101}, {32'b10101010101010101010101010101010, 3'b011}, `__LINE__); // 146: fn=  ADD, a=0x55555555, b=0x55555555, y=0xaaaaaaaa
	test_case({6'b010001, 32'b00000000000000000000000000000000, 32'b00000000000000000000000000000000}, {32'b00000000000000000000000000000000, 3'b100}, `__LINE__); // 147: fn=  SUB, a=0x00000000, b=0x00000000, y=0x00000000
	test_case({6'b010001, 32'b00000000000000000000000000000000, 32'b00000000000000000000000000000001}, {32'b11111111111111111111111111111111, 3'b001}, `__LINE__); // 148: fn=  SUB, a=0x00000000, b=0x00000001, y=0xffffffff
	test_case({6'b010001, 32'b00000000000000000000000000000000, 32'b11111111111111111111111111111111}, {32'b00000000000000000000000000000001, 3'b000}, `__LINE__); // 149: fn=  SUB, a=0x00000000, b=0x-0000001, y=0x00000001
	test_case({6'b010001, 32'b00000000000000000000000000000000, 32'b10101010101010101010101010101010}, {32'b01010101010101010101010101010110, 3'b000}, `__LINE__); // 150: fn=  SUB, a=0x00000000, b=0xaaaaaaaa, y=0x55555556
	test_case({6'b010001, 32'b00000000000000000000000000000000, 32'b01010101010101010101010101010101}, {32'b10101010101010101010101010101011, 3'b001}, `__LINE__); // 151: fn=  SUB, a=0x00000000, b=0x55555555, y=0xaaaaaaab
	test_case({6'b010001, 32'b00000000000000000000000000000001, 32'b00000000000000000000000000000000}, {32'b00000000000000000000000000000001, 3'b000}, `__LINE__); // 152: fn=  SUB, a=0x00000001, b=0x00000000, y=0x00000001
	test_case({6'b010001, 32'b00000000000000000000000000000001, 32'b00000000000000000000000000000001}, {32'b00000000000000000000000000000000, 3'b100}, `__LINE__); // 153: fn=  SUB, a=0x00000001, b=0x00000001, y=0x00000000
	test_case({6'b010001, 32'b00000000000000000000000000000001, 32'b11111111111111111111111111111111}, {32'b00000000000000000000000000000010, 3'b000}, `__LINE__); // 154: fn=  SUB, a=0x00000001, b=0x-0000001, y=0x00000002
	test_case({6'b010001, 32'b00000000000000000000000000000001, 32'b10101010101010101010101010101010}, {32'b01010101010101010101010101010111, 3'b000}, `__LINE__); // 155: fn=  SUB, a=0x00000001, b=0xaaaaaaaa, y=0x55555557
	test_case({6'b010001, 32'b00000000000000000000000000000001, 32'b01010101010101010101010101010101}, {32'b10101010101010101010101010101100, 3'b001}, `__LINE__); // 156: fn=  SUB, a=0x00000001, b=0x55555555, y=0xaaaaaaac
	test_case({6'b010001, 32'b11111111111111111111111111111111, 32'b00000000000000000000000000000000}, {32'b11111111111111111111111111111111, 3'b001}, `__LINE__); // 157: fn=  SUB, a=0x-0000001, b=0x00000000, y=0xffffffff
	test_case({6'b010001, 32'b11111111111111111111111111111111, 32'b00000000000000000000000000000001}, {32'b11111111111111111111111111111110, 3'b001}, `__LINE__); // 158: fn=  SUB, a=0x-0000001, b=0x00000001, y=0xfffffffe
	test_case({6'b010001, 32'b11111111111111111111111111111111, 32'b11111111111111111111111111111111}, {32'b00000000000000000000000000000000, 3'b100}, `__LINE__); // 159: fn=  SUB, a=0x-0000001, b=0x-0000001, y=0x00000000
	test_case({6'b010001, 32'b11111111111111111111111111111111, 32'b10101010101010101010101010101010}, {32'b01010101010101010101010101010101, 3'b000}, `__LINE__); // 160: fn=  SUB, a=0x-0000001, b=0xaaaaaaaa, y=0x55555555
	test_case({6'b010001, 32'b11111111111111111111111111111111, 32'b01010101010101010101010101010101}, {32'b10101010101010101010101010101010, 3'b001}, `__LINE__); // 161: fn=  SUB, a=0x-0000001, b=0x55555555, y=0xaaaaaaaa
	test_case({6'b010001, 32'b10101010101010101010101010101010, 32'b00000000000000000000000000000000}, {32'b10101010101010101010101010101010, 3'b001}, `__LINE__); // 162: fn=  SUB, a=0xaaaaaaaa, b=0x00000000, y=0xaaaaaaaa
	test_case({6'b010001, 32'b10101010101010101010101010101010, 32'b00000000000000000000000000000001}, {32'b10101010101010101010101010101001, 3'b001}, `__LINE__); // 163: fn=  SUB, a=0xaaaaaaaa, b=0x00000001, y=0xaaaaaaa9
	test_case({6'b010001, 32'b10101010101010101010101010101010, 32'b11111111111111111111111111111111}, {32'b10101010101010101010101010101011, 3'b001}, `__LINE__); // 164: fn=  SUB, a=0xaaaaaaaa, b=0x-0000001, y=0xaaaaaaab
	test_case({6'b010001, 32'b10101010101010101010101010101010, 32'b10101010101010101010101010101010}, {32'b00000000000000000000000000000000, 3'b100}, `__LINE__); // 165: fn=  SUB, a=0xaaaaaaaa, b=0xaaaaaaaa, y=0x00000000
	test_case({6'b010001, 32'b10101010101010101010101010101010, 32'b01010101010101010101010101010101}, {32'b01010101010101010101010101010101, 3'b010}, `__LINE__); // 166: fn=  SUB, a=0xaaaaaaaa, b=0x55555555, y=0x55555555
	test_case({6'b010001, 32'b01010101010101010101010101010101, 32'b00000000000000000000000000000000}, {32'b01010101010101010101010101010101, 3'b000}, `__LINE__); // 167: fn=  SUB, a=0x55555555, b=0x00000000, y=0x55555555
	test_case({6'b010001, 32'b01010101010101010101010101010101, 32'b00000000000000000000000000000001}, {32'b01010101010101010101010101010100, 3'b000}, `__LINE__); // 168: fn=  SUB, a=0x55555555, b=0x00000001, y=0x55555554
	test_case({6'b010001, 32'b01010101010101010101010101010101, 32'b11111111111111111111111111111111}, {32'b01010101010101010101010101010110, 3'b000}, `__LINE__); // 169: fn=  SUB, a=0x55555555, b=0x-0000001, y=0x55555556
	test_case({6'b010001, 32'b01010101010101010101010101010101, 32'b10101010101010101010101010101010}, {32'b10101010101010101010101010101011, 3'b011}, `__LINE__); // 170: fn=  SUB, a=0x55555555, b=0xaaaaaaaa, y=0xaaaaaaab
	test_case({6'b010001, 32'b01010101010101010101010101010101, 32'b01010101010101010101010101010101}, {32'b00000000000000000000000000000000, 3'b100}, `__LINE__); // 171: fn=  SUB, a=0x55555555, b=0x55555555, y=0x00000000
	test_case({6'b000011, 32'b00000000000000000000000000000101, 32'b11011110101011011011111011101111}, {32'b00000000000000000000000000000000, 3'b000}, `__LINE__); // 172: fn=CMPEQ, a=0x00000005, b=0xdeadbeef, y=0x00000000
	test_case({6'b000101, 32'b00000000000000000000000000000101, 32'b11011110101011011011111011101111}, {32'b00000000000000000000000000000000, 3'b000}, `__LINE__); // 173: fn=CMPLT, a=0x00000005, b=0xdeadbeef, y=0x00000000
	test_case({6'b000111, 32'b00000000000000000000000000000101, 32'b11011110101011011011111011101111}, {32'b00000000000000000000000000000000, 3'b000}, `__LINE__); // 174: fn=CMPLE, a=0x00000005, b=0xdeadbeef, y=0x00000000
	test_case({6'b000011, 32'b00010010001101000101011001111000, 32'b00010010001101000101011001111000}, {32'b00000000000000000000000000000001, 3'b100}, `__LINE__); // 175: fn=CMPEQ, a=0x12345678, b=0x12345678, y=0x00000001
	test_case({6'b000101, 32'b00010010001101000101011001111000, 32'b00010010001101000101011001111000}, {32'b00000000000000000000000000000000, 3'b100}, `__LINE__); // 176: fn=CMPLT, a=0x12345678, b=0x12345678, y=0x00000000
	test_case({6'b000111, 32'b00010010001101000101011001111000, 32'b00010010001101000101011001111000}, {32'b00000000000000000000000000000001, 3'b100}, `__LINE__); // 177: fn=CMPLE, a=0x12345678, b=0x12345678, y=0x00000001
	test_case({6'b000011, 32'b10000000000000000000000000000000, 32'b00000000000000000000000000000001}, {32'b00000000000000000000000000000000, 3'b010}, `__LINE__); // 178: fn=CMPEQ, a=0x80000000, b=0x00000001, y=0x00000000
	test_case({6'b000101, 32'b10000000000000000000000000000000, 32'b00000000000000000000000000000001}, {32'b00000000000000000000000000000001, 3'b010}, `__LINE__); // 179: fn=CMPLT, a=0x80000000, b=0x00000001, y=0x00000001
	test_case({6'b000111, 32'b10000000000000000000000000000000, 32'b00000000000000000000000000000001}, {32'b00000000000000000000000000000001, 3'b010}, `__LINE__); // 180: fn=CMPLE, a=0x80000000, b=0x00000001, y=0x00000001
	test_case({6'b000011, 32'b11011110101011011011111011101111, 32'b00000000000000000000000000000101}, {32'b00000000000000000000000000000000, 3'b001}, `__LINE__); // 181: fn=CMPEQ, a=0xdeadbeef, b=0x00000005, y=0x00000000
	test_case({6'b000101, 32'b11011110101011011011111011101111, 32'b00000000000000000000000000000101}, {32'b00000000000000000000000000000001, 3'b001}, `__LINE__); // 182: fn=CMPLT, a=0xdeadbeef, b=0x00000005, y=0x00000001
	test_case({6'b000111, 32'b11011110101011011011111011101111, 32'b00000000000000000000000000000101}, {32'b00000000000000000000000000000001, 3'b001}, `__LINE__); // 183: fn=CMPLE, a=0xdeadbeef, b=0x00000005, y=0x00000001
	test_case({6'b000011, 32'b01111111111111111111111111111111, 32'b11111111111111111111111111111111}, {32'b00000000000000000000000000000000, 3'b011}, `__LINE__); // 184: fn=CMPEQ, a=0x7fffffff, b=0xffffffff, y=0x00000000
	test_case({6'b000101, 32'b01111111111111111111111111111111, 32'b11111111111111111111111111111111}, {32'b00000000000000000000000000000000, 3'b011}, `__LINE__); // 185: fn=CMPLT, a=0x7fffffff, b=0xffffffff, y=0x00000000
	test_case({6'b000111, 32'b01111111111111111111111111111111, 32'b11111111111111111111111111111111}, {32'b00000000000000000000000000000000, 3'b011}, `__LINE__); // 186: fn=CMPLE, a=0x7fffffff, b=0xffffffff, y=0x00000000
	$display("");
	if (dut_error != 0) begin
		$display("ERROR: %d test cases failed", dut_error);
		$finish_and_return(1);
	end
	$display("PASS:  all test cases passed");
	$display("");
    $finish;
end


beta_alu dut (
	.a(a),
	.b(b),
    .fn(fn),
    .y(y)
);

endmodule
