// Verilog HDL NetList 
//   timeStamp 2005 7 27 16 43 10 
//   author "Avanti Corporation."
//   program "A2Hdl" 
//   design library: cell
//   cell name     : cell.CEL (version 1)
module SDFFSRX2 ( CK , D , Q , QN , RN , SE , SI , SN );
    input CK ;
    input D ;
    output Q ;
    output QN ;
    input RN ;
    input SE ;
    input SI ;
    input SN ;
endmodule 
module SDFFSRX4 ( CK , D , Q , QN , RN , SE , SI , SN );
    input CK ;
    input D ;
    output Q ;
    output QN ;
    input RN ;
    input SE ;
    input SI ;
    input SN ;
endmodule 
module SDFFSRXL ( CK , D , Q , QN , RN , SE , SI , SN );
    input CK ;
    input D ;
    output Q ;
    output QN ;
    input RN ;
    input SE ;
    input SI ;
    input SN ;
endmodule 
module SDFFSX1 ( CK , D , Q , QN , SE , SI , SN );
    input CK ;
    input D ;
    output Q ;
    output QN ;
    input SE ;
    input SI ;
    input SN ;
endmodule 
module SDFFSX2 ( CK , D , Q , QN , SE , SI , SN );
    input CK ;
    input D ;
    output Q ;
    output QN ;
    input SE ;
    input SI ;
    input SN ;
endmodule 
module SDFFSX4 ( CK , D , Q , QN , SE , SI , SN );
    input CK ;
    input D ;
    output Q ;
    output QN ;
    input SE ;
    input SI ;
    input SN ;
endmodule 
module SDFFSXL ( CK , D , Q , QN , SE , SI , SN );
    input CK ;
    input D ;
    output Q ;
    output QN ;
    input SE ;
    input SI ;
    input SN ;
endmodule 
module SDFFTRX1 ( CK , D , Q , QN , RN , SE , SI );
    input CK ;
    input D ;
    output Q ;
    output QN ;
    input RN ;
    input SE ;
    input SI ;
endmodule 
module SDFFTRX2 ( CK , D , Q , QN , RN , SE , SI );
    input CK ;
    input D ;
    output Q ;
    output QN ;
    input RN ;
    input SE ;
    input SI ;
endmodule 
module SDFFTRX4 ( CK , D , Q , QN , RN , SE , SI );
    input CK ;
    input D ;
    output Q ;
    output QN ;
    input RN ;
    input SE ;
    input SI ;
endmodule 
module SDFFTRXL ( CK , D , Q , QN , RN , SE , SI );
    input CK ;
    input D ;
    output Q ;
    output QN ;
    input RN ;
    input SE ;
    input SI ;
endmodule 
module SDFFX1 ( CK , D , Q , QN , SE , SI );
    input CK ;
    input D ;
    output Q ;
    output QN ;
    input SE ;
    input SI ;
endmodule 
module SDFFX2 ( CK , D , Q , QN , SE , SI );
    input CK ;
    input D ;
    output Q ;
    output QN ;
    input SE ;
    input SI ;
endmodule 
module SMDFFHQX4 ( CK , D0 , D1 , Q , S0 , SE , SI );
    input CK ;
    input D0 ;
    input D1 ;
    output Q ;
    input S0 ;
    input SE ;
    input SI ;
endmodule 
module SMDFFHQX8 ( CK , D0 , D1 , Q , S0 , SE , SI );
    input CK ;
    input D0 ;
    input D1 ;
    output Q ;
    input S0 ;
    input SE ;
    input SI ;
endmodule 
module TBUFX12 ( A , OE , Y );
    input A ;
    input OE ;
    output Y ;
endmodule 
module TBUFX16 ( A , OE , Y );
    input A ;
    input OE ;
    output Y ;
endmodule 
module TBUFX1 ( A , OE , Y );
    input A ;
    input OE ;
    output Y ;
endmodule 
module TBUFX20 ( A , OE , Y );
    input A ;
    input OE ;
    output Y ;
endmodule 
module TBUFX2 ( A , OE , Y );
    input A ;
    input OE ;
    output Y ;
endmodule 
module TBUFX3 ( A , OE , Y );
    input A ;
    input OE ;
    output Y ;
endmodule 
module TBUFX4 ( A , OE , Y );
    input A ;
    input OE ;
    output Y ;
endmodule 
module TBUFX6 ( A , OE , Y );
    input A ;
    input OE ;
    output Y ;
endmodule 
module TBUFX8 ( A , OE , Y );
    input A ;
    input OE ;
    output Y ;
endmodule 
module TBUFXL ( A , OE , Y );
    input A ;
    input OE ;
    output Y ;
endmodule 
module TIEHI ( Y );
    output Y ;
endmodule 
module TIELO ( Y );
    output Y ;
endmodule 
module TLATNCAX12 ( CK , E , ECK );
    input CK ;
    input E ;
    output ECK ;
endmodule 
module TLATNCAX16 ( CK , E , ECK );
    input CK ;
    input E ;
    output ECK ;
endmodule 
module TLATNCAX20 ( CK , E , ECK );
    input CK ;
    input E ;
    output ECK ;
endmodule 
module TLATNCAX2 ( CK , E , ECK );
    input CK ;
    input E ;
    output ECK ;
endmodule 
module TLATNCAX3 ( CK , E , ECK );
    input CK ;
    input E ;
    output ECK ;
endmodule 
module TLATNCAX4 ( CK , E , ECK );
    input CK ;
    input E ;
    output ECK ;
endmodule 
module SDFFSHQX1 ( CK , D , Q , SE , SI , SN );
    input CK ;
    input D ;
    output Q ;
    input SE ;
    input SI ;
    input SN ;
endmodule 
module SDFFSHQX2 ( CK , D , Q , SE , SI , SN );
    input CK ;
    input D ;
    output Q ;
    input SE ;
    input SI ;
    input SN ;
endmodule 
module SDFFSHQX4 ( CK , D , Q , SE , SI , SN );
    input CK ;
    input D ;
    output Q ;
    input SE ;
    input SI ;
    input SN ;
endmodule 
module SDFFSHQX8 ( CK , D , Q , SE , SI , SN );
    input CK ;
    input D ;
    output Q ;
    input SE ;
    input SI ;
    input SN ;
endmodule 
module SDFFSRHQX1 ( CK , D , Q , RN , SE , SI , SN );
    input CK ;
    input D ;
    output Q ;
    input RN ;
    input SE ;
    input SI ;
    input SN ;
endmodule 
module SDFFSRHQX2 ( CK , D , Q , RN , SE , SI , SN );
    input CK ;
    input D ;
    output Q ;
    input RN ;
    input SE ;
    input SI ;
    input SN ;
endmodule 
module SDFFSRHQX4 ( CK , D , Q , RN , SE , SI , SN );
    input CK ;
    input D ;
    output Q ;
    input RN ;
    input SE ;
    input SI ;
    input SN ;
endmodule 
module SDFFSRHQX8 ( CK , D , Q , RN , SE , SI , SN );
    input CK ;
    input D ;
    output Q ;
    input RN ;
    input SE ;
    input SI ;
    input SN ;
endmodule 
module SDFFSRX1 ( CK , D , Q , QN , RN , SE , SI , SN );
    input CK ;
    input D ;
    output Q ;
    output QN ;
    input RN ;
    input SE ;
    input SI ;
    input SN ;
endmodule 
module TLATNTSCAX2 ( CK , E , ECK , SE );
    input CK ;
    input E ;
    output ECK ;
    input SE ;
endmodule 
module TLATNTSCAX3 ( CK , E , ECK , SE );
    input CK ;
    input E ;
    output ECK ;
    input SE ;
endmodule 
module TLATNTSCAX4 ( CK , E , ECK , SE );
    input CK ;
    input E ;
    output ECK ;
    input SE ;
endmodule 
module TLATNTSCAX6 ( CK , E , ECK , SE );
    input CK ;
    input E ;
    output ECK ;
    input SE ;
endmodule 
module TLATNTSCAX8 ( CK , E , ECK , SE );
    input CK ;
    input E ;
    output ECK ;
    input SE ;
endmodule 
module TLATNX1 ( D , GN , Q , QN );
    input D ;
    input GN ;
    output Q ;
    output QN ;
endmodule 
module TLATNX2 ( D , GN , Q , QN );
    input D ;
    input GN ;
    output Q ;
    output QN ;
endmodule 
module TLATNX4 ( D , GN , Q , QN );
    input D ;
    input GN ;
    output Q ;
    output QN ;
endmodule 
module TLATNXL ( D , GN , Q , QN );
    input D ;
    input GN ;
    output Q ;
    output QN ;
endmodule 
module TLATSRX1 ( D , G , Q , QN , RN , SN );
    input D ;
    input G ;
    output Q ;
    output QN ;
    input RN ;
    input SN ;
endmodule 
module TLATSRX2 ( D , G , Q , QN , RN , SN );
    input D ;
    input G ;
    output Q ;
    output QN ;
    input RN ;
    input SN ;
endmodule 
module TLATSRX4 ( D , G , Q , QN , RN , SN );
    input D ;
    input G ;
    output Q ;
    output QN ;
    input RN ;
    input SN ;
endmodule 
module TLATSRXL ( D , G , Q , QN , RN , SN );
    input D ;
    input G ;
    output Q ;
    output QN ;
    input RN ;
    input SN ;
endmodule 
module TLATX1 ( D , G , Q , QN );
    input D ;
    input G ;
    output Q ;
    output QN ;
endmodule 
module TLATX2 ( D , G , Q , QN );
    input D ;
    input G ;
    output Q ;
    output QN ;
endmodule 
module TLATX4 ( D , G , Q , QN );
    input D ;
    input G ;
    output Q ;
    output QN ;
endmodule 
module TLATXL ( D , G , Q , QN );
    input D ;
    input G ;
    output Q ;
    output QN ;
endmodule 
module XNOR2X1 ( A , B , Y );
    input A ;
    input B ;
    output Y ;
endmodule 
module XNOR2X2 ( A , B , Y );
    input A ;
    input B ;
    output Y ;
endmodule 
module XNOR2X4 ( A , B , Y );
    input A ;
    input B ;
    output Y ;
endmodule 
module SEDFFTRX2 ( CK , D , E , Q , QN , RN , SE , SI );
    input CK ;
    input D ;
    input E ;
    output Q ;
    output QN ;
    input RN ;
    input SE ;
    input SI ;
endmodule 
module SEDFFTRX4 ( CK , D , E , Q , QN , RN , SE , SI );
    input CK ;
    input D ;
    input E ;
    output Q ;
    output QN ;
    input RN ;
    input SE ;
    input SI ;
endmodule 
module SEDFFTRXL ( CK , D , E , Q , QN , RN , SE , SI );
    input CK ;
    input D ;
    input E ;
    output Q ;
    output QN ;
    input RN ;
    input SE ;
    input SI ;
endmodule 
module SEDFFX1 ( CK , D , E , Q , QN , SE , SI );
    input CK ;
    input D ;
    input E ;
    output Q ;
    output QN ;
    input SE ;
    input SI ;
endmodule 
module SEDFFX2 ( CK , D , E , Q , QN , SE , SI );
    input CK ;
    input D ;
    input E ;
    output Q ;
    output QN ;
    input SE ;
    input SI ;
endmodule 
module SEDFFX4 ( CK , D , E , Q , QN , SE , SI );
    input CK ;
    input D ;
    input E ;
    output Q ;
    output QN ;
    input SE ;
    input SI ;
endmodule 
module SEDFFXL ( CK , D , E , Q , QN , SE , SI );
    input CK ;
    input D ;
    input E ;
    output Q ;
    output QN ;
    input SE ;
    input SI ;
endmodule 
module SMDFFHQX1 ( CK , D0 , D1 , Q , S0 , SE , SI );
    input CK ;
    input D0 ;
    input D1 ;
    output Q ;
    input S0 ;
    input SE ;
    input SI ;
endmodule 
module SMDFFHQX2 ( CK , D0 , D1 , Q , S0 , SE , SI );
    input CK ;
    input D0 ;
    input D1 ;
    output Q ;
    input S0 ;
    input SE ;
    input SI ;
endmodule 
module OAI22X2 ( A0 , A1 , B0 , B1 , Y );
    input A0 ;
    input A1 ;
    input B0 ;
    input B1 ;
    output Y ;
endmodule 
module OAI22X4 ( A0 , A1 , B0 , B1 , Y );
    input A0 ;
    input A1 ;
    input B0 ;
    input B1 ;
    output Y ;
endmodule 
module OAI22XL ( A0 , A1 , B0 , B1 , Y );
    input A0 ;
    input A1 ;
    input B0 ;
    input B1 ;
    output Y ;
endmodule 
module OAI2BB1X1 ( A0N , A1N , B0 , Y );
    input A0N ;
    input A1N ;
    input B0 ;
    output Y ;
endmodule 
module OAI2BB1X2 ( A0N , A1N , B0 , Y );
    input A0N ;
    input A1N ;
    input B0 ;
    output Y ;
endmodule 
module OAI2BB1X4 ( A0N , A1N , B0 , Y );
    input A0N ;
    input A1N ;
    input B0 ;
    output Y ;
endmodule 
module OAI2BB1XL ( A0N , A1N , B0 , Y );
    input A0N ;
    input A1N ;
    input B0 ;
    output Y ;
endmodule 
module XNOR2XL ( A , B , Y );
    input A ;
    input B ;
    output Y ;
endmodule 
module XNOR3X1 ( A , B , C , Y );
    input A ;
    input B ;
    input C ;
    output Y ;
endmodule 
module XNOR3X2 ( A , B , C , Y );
    input A ;
    input B ;
    input C ;
    output Y ;
endmodule 
module XNOR3X4 ( A , B , C , Y );
    input A ;
    input B ;
    input C ;
    output Y ;
endmodule 
module XNOR3XL ( A , B , C , Y );
    input A ;
    input B ;
    input C ;
    output Y ;
endmodule 
module XOR2X1 ( A , B , Y );
    input A ;
    input B ;
    output Y ;
endmodule 
module XOR2X2 ( A , B , Y );
    input A ;
    input B ;
    output Y ;
endmodule 
module XOR2X4 ( A , B , Y );
    input A ;
    input B ;
    output Y ;
endmodule 
module XOR2XL ( A , B , Y );
    input A ;
    input B ;
    output Y ;
endmodule 
module XOR3X1 ( A , B , C , Y );
    input A ;
    input B ;
    input C ;
    output Y ;
endmodule 
module XOR3X2 ( A , B , C , Y );
    input A ;
    input B ;
    input C ;
    output Y ;
endmodule 
module XOR3X4 ( A , B , C , Y );
    input A ;
    input B ;
    input C ;
    output Y ;
endmodule 
module XOR3XL ( A , B , C , Y );
    input A ;
    input B ;
    input C ;
    output Y ;
endmodule 
module TLATNCAX6 ( CK , E , ECK );
    input CK ;
    input E ;
    output ECK ;
endmodule 
module TLATNCAX8 ( CK , E , ECK );
    input CK ;
    input E ;
    output ECK ;
endmodule 
module TLATNSRX1 ( D , GN , Q , QN , RN , SN );
    input D ;
    input GN ;
    output Q ;
    output QN ;
    input RN ;
    input SN ;
endmodule 
module TLATNSRX2 ( D , GN , Q , QN , RN , SN );
    input D ;
    input GN ;
    output Q ;
    output QN ;
    input RN ;
    input SN ;
endmodule 
module TLATNSRX4 ( D , GN , Q , QN , RN , SN );
    input D ;
    input GN ;
    output Q ;
    output QN ;
    input RN ;
    input SN ;
endmodule 
module TLATNSRXL ( D , GN , Q , QN , RN , SN );
    input D ;
    input GN ;
    output Q ;
    output QN ;
    input RN ;
    input SN ;
endmodule 
module TLATNTSCAX12 ( CK , E , ECK , SE );
    input CK ;
    input E ;
    output ECK ;
    input SE ;
endmodule 
module TLATNTSCAX16 ( CK , E , ECK , SE );
    input CK ;
    input E ;
    output ECK ;
    input SE ;
endmodule 
module TLATNTSCAX20 ( CK , E , ECK , SE );
    input CK ;
    input E ;
    output ECK ;
    input SE ;
endmodule 
module OR3X1 ( A , B , C , Y );
    input A ;
    input B ;
    input C ;
    output Y ;
endmodule 
module OR3X2 ( A , B , C , Y );
    input A ;
    input B ;
    input C ;
    output Y ;
endmodule 
module OR3X4 ( A , B , C , Y );
    input A ;
    input B ;
    input C ;
    output Y ;
endmodule 
module OR3X6 ( A , B , C , Y );
    input A ;
    input B ;
    input C ;
    output Y ;
endmodule 
module OR3X8 ( A , B , C , Y );
    input A ;
    input B ;
    input C ;
    output Y ;
endmodule 
module OR3XL ( A , B , C , Y );
    input A ;
    input B ;
    input C ;
    output Y ;
endmodule 
module OR4X1 ( A , B , C , D , Y );
    input A ;
    input B ;
    input C ;
    input D ;
    output Y ;
endmodule 
module OR4X2 ( A , B , C , D , Y );
    input A ;
    input B ;
    input C ;
    input D ;
    output Y ;
endmodule 
module OA22X1 ( A0 , A1 , B0 , B1 , Y );
    input A0 ;
    input A1 ;
    input B0 ;
    input B1 ;
    output Y ;
endmodule 
module OA22X2 ( A0 , A1 , B0 , B1 , Y );
    input A0 ;
    input A1 ;
    input B0 ;
    input B1 ;
    output Y ;
endmodule 
module OA22X4 ( A0 , A1 , B0 , B1 , Y );
    input A0 ;
    input A1 ;
    input B0 ;
    input B1 ;
    output Y ;
endmodule 
module OA22XL ( A0 , A1 , B0 , B1 , Y );
    input A0 ;
    input A1 ;
    input B0 ;
    input B1 ;
    output Y ;
endmodule 
module OAI211X1 ( A0 , A1 , B0 , C0 , Y );
    input A0 ;
    input A1 ;
    input B0 ;
    input C0 ;
    output Y ;
endmodule 
module OAI211X2 ( A0 , A1 , B0 , C0 , Y );
    input A0 ;
    input A1 ;
    input B0 ;
    input C0 ;
    output Y ;
endmodule 
module OAI211X4 ( A0 , A1 , B0 , C0 , Y );
    input A0 ;
    input A1 ;
    input B0 ;
    input C0 ;
    output Y ;
endmodule 
module OAI211XL ( A0 , A1 , B0 , C0 , Y );
    input A0 ;
    input A1 ;
    input B0 ;
    input C0 ;
    output Y ;
endmodule 
module OAI21X1 ( A0 , A1 , B0 , Y );
    input A0 ;
    input A1 ;
    input B0 ;
    output Y ;
endmodule 
module OAI21X2 ( A0 , A1 , B0 , Y );
    input A0 ;
    input A1 ;
    input B0 ;
    output Y ;
endmodule 
module OAI21X4 ( A0 , A1 , B0 , Y );
    input A0 ;
    input A1 ;
    input B0 ;
    output Y ;
endmodule 
module OAI21XL ( A0 , A1 , B0 , Y );
    input A0 ;
    input A1 ;
    input B0 ;
    output Y ;
endmodule 
module OAI221X1 ( A0 , A1 , B0 , B1 , C0 , Y );
    input A0 ;
    input A1 ;
    input B0 ;
    input B1 ;
    input C0 ;
    output Y ;
endmodule 
module OAI221X2 ( A0 , A1 , B0 , B1 , C0 , Y );
    input A0 ;
    input A1 ;
    input B0 ;
    input B1 ;
    input C0 ;
    output Y ;
endmodule 
module OAI221X4 ( A0 , A1 , B0 , B1 , C0 , Y );
    input A0 ;
    input A1 ;
    input B0 ;
    input B1 ;
    input C0 ;
    output Y ;
endmodule 
module OAI221XL ( A0 , A1 , B0 , B1 , C0 , Y );
    input A0 ;
    input A1 ;
    input B0 ;
    input B1 ;
    input C0 ;
    output Y ;
endmodule 
module OAI222X1 ( A0 , A1 , B0 , B1 , C0 , C1 , Y );
    input A0 ;
    input A1 ;
    input B0 ;
    input B1 ;
    input C0 ;
    input C1 ;
    output Y ;
endmodule 
module OAI222X2 ( A0 , A1 , B0 , B1 , C0 , C1 , Y );
    input A0 ;
    input A1 ;
    input B0 ;
    input B1 ;
    input C0 ;
    input C1 ;
    output Y ;
endmodule 
module OAI222X4 ( A0 , A1 , B0 , B1 , C0 , C1 , Y );
    input A0 ;
    input A1 ;
    input B0 ;
    input B1 ;
    input C0 ;
    input C1 ;
    output Y ;
endmodule 
module OAI222XL ( A0 , A1 , B0 , B1 , C0 , C1 , Y );
    input A0 ;
    input A1 ;
    input B0 ;
    input B1 ;
    input C0 ;
    input C1 ;
    output Y ;
endmodule 
module OAI22X1 ( A0 , A1 , B0 , B1 , Y );
    input A0 ;
    input A1 ;
    input B0 ;
    input B1 ;
    output Y ;
endmodule 
module SDFFRHQX1 ( CK , D , Q , RN , SE , SI );
    input CK ;
    input D ;
    output Q ;
    input RN ;
    input SE ;
    input SI ;
endmodule 
module SDFFRHQX2 ( CK , D , Q , RN , SE , SI );
    input CK ;
    input D ;
    output Q ;
    input RN ;
    input SE ;
    input SI ;
endmodule 
module SDFFRHQX4 ( CK , D , Q , RN , SE , SI );
    input CK ;
    input D ;
    output Q ;
    input RN ;
    input SE ;
    input SI ;
endmodule 
module SDFFRHQX8 ( CK , D , Q , RN , SE , SI );
    input CK ;
    input D ;
    output Q ;
    input RN ;
    input SE ;
    input SI ;
endmodule 
module SDFFRX1 ( CK , D , Q , QN , RN , SE , SI );
    input CK ;
    input D ;
    output Q ;
    output QN ;
    input RN ;
    input SE ;
    input SI ;
endmodule 
module SDFFRX2 ( CK , D , Q , QN , RN , SE , SI );
    input CK ;
    input D ;
    output Q ;
    output QN ;
    input RN ;
    input SE ;
    input SI ;
endmodule 
module SDFFRX4 ( CK , D , Q , QN , RN , SE , SI );
    input CK ;
    input D ;
    output Q ;
    output QN ;
    input RN ;
    input SE ;
    input SI ;
endmodule 
module SDFFRXL ( CK , D , Q , QN , RN , SE , SI );
    input CK ;
    input D ;
    output Q ;
    output QN ;
    input RN ;
    input SE ;
    input SI ;
endmodule 
module OAI2BB2X2 ( A0N , A1N , B0 , B1 , Y );
    input A0N ;
    input A1N ;
    input B0 ;
    input B1 ;
    output Y ;
endmodule 
module OAI2BB2X4 ( A0N , A1N , B0 , B1 , Y );
    input A0N ;
    input A1N ;
    input B0 ;
    input B1 ;
    output Y ;
endmodule 
module OAI2BB2XL ( A0N , A1N , B0 , B1 , Y );
    input A0N ;
    input A1N ;
    input B0 ;
    input B1 ;
    output Y ;
endmodule 
module OAI31X1 ( A0 , A1 , A2 , B0 , Y );
    input A0 ;
    input A1 ;
    input A2 ;
    input B0 ;
    output Y ;
endmodule 
module OAI31X2 ( A0 , A1 , A2 , B0 , Y );
    input A0 ;
    input A1 ;
    input A2 ;
    input B0 ;
    output Y ;
endmodule 
module OAI31X4 ( A0 , A1 , A2 , B0 , Y );
    input A0 ;
    input A1 ;
    input A2 ;
    input B0 ;
    output Y ;
endmodule 
module OAI31XL ( A0 , A1 , A2 , B0 , Y );
    input A0 ;
    input A1 ;
    input A2 ;
    input B0 ;
    output Y ;
endmodule 
module OAI32X1 ( A0 , A1 , A2 , B0 , B1 , Y );
    input A0 ;
    input A1 ;
    input A2 ;
    input B0 ;
    input B1 ;
    output Y ;
endmodule 
module OAI32X2 ( A0 , A1 , A2 , B0 , B1 , Y );
    input A0 ;
    input A1 ;
    input A2 ;
    input B0 ;
    input B1 ;
    output Y ;
endmodule 
module OAI32X4 ( A0 , A1 , A2 , B0 , B1 , Y );
    input A0 ;
    input A1 ;
    input A2 ;
    input B0 ;
    input B1 ;
    output Y ;
endmodule 
module OAI32XL ( A0 , A1 , A2 , B0 , B1 , Y );
    input A0 ;
    input A1 ;
    input A2 ;
    input B0 ;
    input B1 ;
    output Y ;
endmodule 
module OAI33X1 ( A0 , A1 , A2 , B0 , B1 , B2 , Y );
    input A0 ;
    input A1 ;
    input A2 ;
    input B0 ;
    input B1 ;
    input B2 ;
    output Y ;
endmodule 
module OAI33X2 ( A0 , A1 , A2 , B0 , B1 , B2 , Y );
    input A0 ;
    input A1 ;
    input A2 ;
    input B0 ;
    input B1 ;
    input B2 ;
    output Y ;
endmodule 
module OAI33X4 ( A0 , A1 , A2 , B0 , B1 , B2 , Y );
    input A0 ;
    input A1 ;
    input A2 ;
    input B0 ;
    input B1 ;
    input B2 ;
    output Y ;
endmodule 
module OAI33XL ( A0 , A1 , A2 , B0 , B1 , B2 , Y );
    input A0 ;
    input A1 ;
    input A2 ;
    input B0 ;
    input B1 ;
    input B2 ;
    output Y ;
endmodule 
module OR2X1 ( A , B , Y );
    input A ;
    input B ;
    output Y ;
endmodule 
module OR2X2 ( A , B , Y );
    input A ;
    input B ;
    output Y ;
endmodule 
module OR2X4 ( A , B , Y );
    input A ;
    input B ;
    output Y ;
endmodule 
module OR2X6 ( A , B , Y );
    input A ;
    input B ;
    output Y ;
endmodule 
module OR2X8 ( A , B , Y );
    input A ;
    input B ;
    output Y ;
endmodule 
module OR2XL ( A , B , Y );
    input A ;
    input B ;
    output Y ;
endmodule 
module INVX1 ( A , Y );
    input A ;
    output Y ;
endmodule 
module SDFFX4 ( CK , D , Q , QN , SE , SI );
    input CK ;
    input D ;
    output Q ;
    output QN ;
    input SE ;
    input SI ;
endmodule 
module SDFFXL ( CK , D , Q , QN , SE , SI );
    input CK ;
    input D ;
    output Q ;
    output QN ;
    input SE ;
    input SI ;
endmodule 
module SEDFFHQX1 ( CK , D , E , Q , SE , SI );
    input CK ;
    input D ;
    input E ;
    output Q ;
    input SE ;
    input SI ;
endmodule 
module SEDFFHQX2 ( CK , D , E , Q , SE , SI );
    input CK ;
    input D ;
    input E ;
    output Q ;
    input SE ;
    input SI ;
endmodule 
module SEDFFHQX4 ( CK , D , E , Q , SE , SI );
    input CK ;
    input D ;
    input E ;
    output Q ;
    input SE ;
    input SI ;
endmodule 
module SEDFFHQX8 ( CK , D , E , Q , SE , SI );
    input CK ;
    input D ;
    input E ;
    output Q ;
    input SE ;
    input SI ;
endmodule 
module SEDFFTRX1 ( CK , D , E , Q , QN , RN , SE , SI );
    input CK ;
    input D ;
    input E ;
    output Q ;
    output QN ;
    input RN ;
    input SE ;
    input SI ;
endmodule 
module OR4X4 ( A , B , C , D , Y );
    input A ;
    input B ;
    input C ;
    input D ;
    output Y ;
endmodule 
module OR4X6 ( A , B , C , D , Y );
    input A ;
    input B ;
    input C ;
    input D ;
    output Y ;
endmodule 
module OR4X8 ( A , B , C , D , Y );
    input A ;
    input B ;
    input C ;
    input D ;
    output Y ;
endmodule 
module OR4XL ( A , B , C , D , Y );
    input A ;
    input B ;
    input C ;
    input D ;
    output Y ;
endmodule 
module RF1R1WX1 ( RB , RW , RWN , WB , WW );
    output RB ;
    input RW ;
    input RWN ;
    input WB ;
    input WW ;
endmodule 
module RF2R1WX1 ( R1B , R1W , R2B , R2W , WB , WW );
    output R1B ;
    input R1W ;
    output R2B ;
    input R2W ;
    input WB ;
    input WW ;
endmodule 
module RFRDX1 ( BRB , RB );
    output BRB ;
    input RB ;
endmodule 
module RFRDX2 ( BRB , RB );
    output BRB ;
    input RB ;
endmodule 
module RFRDX4 ( BRB , RB );
    output BRB ;
    input RB ;
endmodule 
module SDFFHQX1 ( CK , D , Q , SE , SI );
    input CK ;
    input D ;
    output Q ;
    input SE ;
    input SI ;
endmodule 
module SDFFHQX2 ( CK , D , Q , SE , SI );
    input CK ;
    input D ;
    output Q ;
    input SE ;
    input SI ;
endmodule 
module SDFFHQX4 ( CK , D , Q , SE , SI );
    input CK ;
    input D ;
    output Q ;
    input SE ;
    input SI ;
endmodule 
module SDFFHQX8 ( CK , D , Q , SE , SI );
    input CK ;
    input D ;
    output Q ;
    input SE ;
    input SI ;
endmodule 
module SDFFNSRX1 ( CKN , D , Q , QN , RN , SE , SI , SN );
    input CKN ;
    input D ;
    output Q ;
    output QN ;
    input RN ;
    input SE ;
    input SI ;
    input SN ;
endmodule 
module SDFFNSRX2 ( CKN , D , Q , QN , RN , SE , SI , SN );
    input CKN ;
    input D ;
    output Q ;
    output QN ;
    input RN ;
    input SE ;
    input SI ;
    input SN ;
endmodule 
module SDFFNSRX4 ( CKN , D , Q , QN , RN , SE , SI , SN );
    input CKN ;
    input D ;
    output Q ;
    output QN ;
    input RN ;
    input SE ;
    input SI ;
    input SN ;
endmodule 
module SDFFNSRXL ( CKN , D , Q , QN , RN , SE , SI , SN );
    input CKN ;
    input D ;
    output Q ;
    output QN ;
    input RN ;
    input SE ;
    input SI ;
    input SN ;
endmodule 
module SDFFQX1 ( CK , D , Q , SE , SI );
    input CK ;
    input D ;
    output Q ;
    input SE ;
    input SI ;
endmodule 
module SDFFQX2 ( CK , D , Q , SE , SI );
    input CK ;
    input D ;
    output Q ;
    input SE ;
    input SI ;
endmodule 
module SDFFQX4 ( CK , D , Q , SE , SI );
    input CK ;
    input D ;
    output Q ;
    input SE ;
    input SI ;
endmodule 
module SDFFQXL ( CK , D , Q , SE , SI );
    input CK ;
    input D ;
    output Q ;
    input SE ;
    input SI ;
endmodule 
module MXI2X6 ( A , B , S0 , Y );
    input A ;
    input B ;
    input S0 ;
    output Y ;
endmodule 
module MXI2X8 ( A , B , S0 , Y );
    input A ;
    input B ;
    input S0 ;
    output Y ;
endmodule 
module MXI2XL ( A , B , S0 , Y );
    input A ;
    input B ;
    input S0 ;
    output Y ;
endmodule 
module MXI3X1 ( A , B , C , S0 , S1 , Y );
    input A ;
    input B ;
    input C ;
    input S0 ;
    input S1 ;
    output Y ;
endmodule 
module MXI3X2 ( A , B , C , S0 , S1 , Y );
    input A ;
    input B ;
    input C ;
    input S0 ;
    input S1 ;
    output Y ;
endmodule 
module MXI3X4 ( A , B , C , S0 , S1 , Y );
    input A ;
    input B ;
    input C ;
    input S0 ;
    input S1 ;
    output Y ;
endmodule 
module MXI3XL ( A , B , C , S0 , S1 , Y );
    input A ;
    input B ;
    input C ;
    input S0 ;
    input S1 ;
    output Y ;
endmodule 
module MXI4X1 ( A , B , C , D , S0 , S1 , Y );
    input A ;
    input B ;
    input C ;
    input D ;
    input S0 ;
    input S1 ;
    output Y ;
endmodule 
module MXI4X2 ( A , B , C , D , S0 , S1 , Y );
    input A ;
    input B ;
    input C ;
    input D ;
    input S0 ;
    input S1 ;
    output Y ;
endmodule 
module MXI4X4 ( A , B , C , D , S0 , S1 , Y );
    input A ;
    input B ;
    input C ;
    input D ;
    input S0 ;
    input S1 ;
    output Y ;
endmodule 
module MXI4XL ( A , B , C , D , S0 , S1 , Y );
    input A ;
    input B ;
    input C ;
    input D ;
    input S0 ;
    input S1 ;
    output Y ;
endmodule 
module NAND2BX1 ( AN , B , Y );
    input AN ;
    input B ;
    output Y ;
endmodule 
module NAND2BX2 ( AN , B , Y );
    input AN ;
    input B ;
    output Y ;
endmodule 
module NAND2BX4 ( AN , B , Y );
    input AN ;
    input B ;
    output Y ;
endmodule 
module NAND2BXL ( AN , B , Y );
    input AN ;
    input B ;
    output Y ;
endmodule 
module NAND2X1 ( A , B , Y );
    input A ;
    input B ;
    output Y ;
endmodule 
module NAND2X2 ( A , B , Y );
    input A ;
    input B ;
    output Y ;
endmodule 
module NAND2X4 ( A , B , Y );
    input A ;
    input B ;
    output Y ;
endmodule 
module NAND2X6 ( A , B , Y );
    input A ;
    input B ;
    output Y ;
endmodule 
module NAND2X8 ( A , B , Y );
    input A ;
    input B ;
    output Y ;
endmodule 
module NAND2XL ( A , B , Y );
    input A ;
    input B ;
    output Y ;
endmodule 
module NAND3BX1 ( AN , B , C , Y );
    input AN ;
    input B ;
    input C ;
    output Y ;
endmodule 
module NAND3BX2 ( AN , B , C , Y );
    input AN ;
    input B ;
    input C ;
    output Y ;
endmodule 
module NAND3BX4 ( AN , B , C , Y );
    input AN ;
    input B ;
    input C ;
    output Y ;
endmodule 
module NAND3BXL ( AN , B , C , Y );
    input AN ;
    input B ;
    input C ;
    output Y ;
endmodule 
module FILL8 ();
endmodule 
module HOLDX1 ( Y );
    inout Y ;
endmodule 
module INVX12 ( A , Y );
    input A ;
    output Y ;
endmodule 
module INVX16 ( A , Y );
    input A ;
    output Y ;
endmodule 
module NAND3X8 ( A , B , C , Y );
    input A ;
    input B ;
    input C ;
    output Y ;
endmodule 
module NAND3XL ( A , B , C , Y );
    input A ;
    input B ;
    input C ;
    output Y ;
endmodule 
module NAND4BBX1 ( AN , BN , C , D , Y );
    input AN ;
    input BN ;
    input C ;
    input D ;
    output Y ;
endmodule 
module NAND4BBX2 ( AN , BN , C , D , Y );
    input AN ;
    input BN ;
    input C ;
    input D ;
    output Y ;
endmodule 
module NAND4BBX4 ( AN , BN , C , D , Y );
    input AN ;
    input BN ;
    input C ;
    input D ;
    output Y ;
endmodule 
module NAND4BBXL ( AN , BN , C , D , Y );
    input AN ;
    input BN ;
    input C ;
    input D ;
    output Y ;
endmodule 
module NAND4BX1 ( AN , B , C , D , Y );
    input AN ;
    input B ;
    input C ;
    input D ;
    output Y ;
endmodule 
module NAND4BX2 ( AN , B , C , D , Y );
    input AN ;
    input B ;
    input C ;
    input D ;
    output Y ;
endmodule 
module NAND4BX4 ( AN , B , C , D , Y );
    input AN ;
    input B ;
    input C ;
    input D ;
    output Y ;
endmodule 
module NAND4BXL ( AN , B , C , D , Y );
    input AN ;
    input B ;
    input C ;
    input D ;
    output Y ;
endmodule 
module NAND4X1 ( A , B , C , D , Y );
    input A ;
    input B ;
    input C ;
    input D ;
    output Y ;
endmodule 
module NAND4X2 ( A , B , C , D , Y );
    input A ;
    input B ;
    input C ;
    input D ;
    output Y ;
endmodule 
module NAND4X4 ( A , B , C , D , Y );
    input A ;
    input B ;
    input C ;
    input D ;
    output Y ;
endmodule 
module NAND4X6 ( A , B , C , D , Y );
    input A ;
    input B ;
    input C ;
    input D ;
    output Y ;
endmodule 
module NAND4X8 ( A , B , C , D , Y );
    input A ;
    input B ;
    input C ;
    input D ;
    output Y ;
endmodule 
module NAND4XL ( A , B , C , D , Y );
    input A ;
    input B ;
    input C ;
    input D ;
    output Y ;
endmodule 
module NOR2BX1 ( AN , B , Y );
    input AN ;
    input B ;
    output Y ;
endmodule 
module NOR2BX2 ( AN , B , Y );
    input AN ;
    input B ;
    output Y ;
endmodule 
module NOR2BX4 ( AN , B , Y );
    input AN ;
    input B ;
    output Y ;
endmodule 
module NOR2BXL ( AN , B , Y );
    input AN ;
    input B ;
    output Y ;
endmodule 
module NOR2X1 ( A , B , Y );
    input A ;
    input B ;
    output Y ;
endmodule 
module NOR2X2 ( A , B , Y );
    input A ;
    input B ;
    output Y ;
endmodule 
module NOR2X4 ( A , B , Y );
    input A ;
    input B ;
    output Y ;
endmodule 
module NOR2X6 ( A , B , Y );
    input A ;
    input B ;
    output Y ;
endmodule 
module NOR2X8 ( A , B , Y );
    input A ;
    input B ;
    output Y ;
endmodule 
module MX4XL ( A , B , C , D , S0 , S1 , Y );
    input A ;
    input B ;
    input C ;
    input D ;
    input S0 ;
    input S1 ;
    output Y ;
endmodule 
module MXI2X1 ( A , B , S0 , Y );
    input A ;
    input B ;
    input S0 ;
    output Y ;
endmodule 
module MXI2X2 ( A , B , S0 , Y );
    input A ;
    input B ;
    input S0 ;
    output Y ;
endmodule 
module MXI2X4 ( A , B , S0 , Y );
    input A ;
    input B ;
    input S0 ;
    output Y ;
endmodule 
module NOR3BXL ( AN , B , C , Y );
    input AN ;
    input B ;
    input C ;
    output Y ;
endmodule 
module NOR3X1 ( A , B , C , Y );
    input A ;
    input B ;
    input C ;
    output Y ;
endmodule 
module NOR3X2 ( A , B , C , Y );
    input A ;
    input B ;
    input C ;
    output Y ;
endmodule 
module NOR3X4 ( A , B , C , Y );
    input A ;
    input B ;
    input C ;
    output Y ;
endmodule 
module NOR3X6 ( A , B , C , Y );
    input A ;
    input B ;
    input C ;
    output Y ;
endmodule 
module NOR3X8 ( A , B , C , Y );
    input A ;
    input B ;
    input C ;
    output Y ;
endmodule 
module NOR3XL ( A , B , C , Y );
    input A ;
    input B ;
    input C ;
    output Y ;
endmodule 
module NOR4BBX1 ( AN , BN , C , D , Y );
    input AN ;
    input BN ;
    input C ;
    input D ;
    output Y ;
endmodule 
module NOR4BBX2 ( AN , BN , C , D , Y );
    input AN ;
    input BN ;
    input C ;
    input D ;
    output Y ;
endmodule 
module NOR4BBX4 ( AN , BN , C , D , Y );
    input AN ;
    input BN ;
    input C ;
    input D ;
    output Y ;
endmodule 
module NOR4BBXL ( AN , BN , C , D , Y );
    input AN ;
    input BN ;
    input C ;
    input D ;
    output Y ;
endmodule 
module NOR4BX1 ( AN , B , C , D , Y );
    input AN ;
    input B ;
    input C ;
    input D ;
    output Y ;
endmodule 
module NOR4BX2 ( AN , B , C , D , Y );
    input AN ;
    input B ;
    input C ;
    input D ;
    output Y ;
endmodule 
module NOR4BX4 ( AN , B , C , D , Y );
    input AN ;
    input B ;
    input C ;
    input D ;
    output Y ;
endmodule 
module NOR4BXL ( AN , B , C , D , Y );
    input AN ;
    input B ;
    input C ;
    input D ;
    output Y ;
endmodule 
module NOR4X1 ( A , B , C , D , Y );
    input A ;
    input B ;
    input C ;
    input D ;
    output Y ;
endmodule 
module NOR4X2 ( A , B , C , D , Y );
    input A ;
    input B ;
    input C ;
    input D ;
    output Y ;
endmodule 
module NOR4X4 ( A , B , C , D , Y );
    input A ;
    input B ;
    input C ;
    input D ;
    output Y ;
endmodule 
module NOR4X6 ( A , B , C , D , Y );
    input A ;
    input B ;
    input C ;
    input D ;
    output Y ;
endmodule 
module NOR4X8 ( A , B , C , D , Y );
    input A ;
    input B ;
    input C ;
    input D ;
    output Y ;
endmodule 
module NOR4XL ( A , B , C , D , Y );
    input A ;
    input B ;
    input C ;
    input D ;
    output Y ;
endmodule 
module OA21X1 ( A0 , A1 , B0 , Y );
    input A0 ;
    input A1 ;
    input B0 ;
    output Y ;
endmodule 
module OA21X2 ( A0 , A1 , B0 , Y );
    input A0 ;
    input A1 ;
    input B0 ;
    output Y ;
endmodule 
module OA21X4 ( A0 , A1 , B0 , Y );
    input A0 ;
    input A1 ;
    input B0 ;
    output Y ;
endmodule 
module OA21XL ( A0 , A1 , B0 , Y );
    input A0 ;
    input A1 ;
    input B0 ;
    output Y ;
endmodule 
module NAND3X1 ( A , B , C , Y );
    input A ;
    input B ;
    input C ;
    output Y ;
endmodule 
module NAND3X2 ( A , B , C , Y );
    input A ;
    input B ;
    input C ;
    output Y ;
endmodule 
module NAND3X4 ( A , B , C , Y );
    input A ;
    input B ;
    input C ;
    output Y ;
endmodule 
module NAND3X6 ( A , B , C , Y );
    input A ;
    input B ;
    input C ;
    output Y ;
endmodule 
module DFFSRX1 ( CK , D , Q , QN , RN , SN );
    input CK ;
    input D ;
    output Q ;
    output QN ;
    input RN ;
    input SN ;
endmodule 
module DFFSRX2 ( CK , D , Q , QN , RN , SN );
    input CK ;
    input D ;
    output Q ;
    output QN ;
    input RN ;
    input SN ;
endmodule 
module DFFSRX4 ( CK , D , Q , QN , RN , SN );
    input CK ;
    input D ;
    output Q ;
    output QN ;
    input RN ;
    input SN ;
endmodule 
module DFFSRXL ( CK , D , Q , QN , RN , SN );
    input CK ;
    input D ;
    output Q ;
    output QN ;
    input RN ;
    input SN ;
endmodule 
module DFFSX1 ( CK , D , Q , QN , SN );
    input CK ;
    input D ;
    output Q ;
    output QN ;
    input SN ;
endmodule 
module DFFSX2 ( CK , D , Q , QN , SN );
    input CK ;
    input D ;
    output Q ;
    output QN ;
    input SN ;
endmodule 
module DFFSX4 ( CK , D , Q , QN , SN );
    input CK ;
    input D ;
    output Q ;
    output QN ;
    input SN ;
endmodule 
module DFFSXL ( CK , D , Q , QN , SN );
    input CK ;
    input D ;
    output Q ;
    output QN ;
    input SN ;
endmodule 
module DFFTRX1 ( CK , D , Q , QN , RN );
    input CK ;
    input D ;
    output Q ;
    output QN ;
    input RN ;
endmodule 
module DFFTRX2 ( CK , D , Q , QN , RN );
    input CK ;
    input D ;
    output Q ;
    output QN ;
    input RN ;
endmodule 
module DFFTRX4 ( CK , D , Q , QN , RN );
    input CK ;
    input D ;
    output Q ;
    output QN ;
    input RN ;
endmodule 
module DFFTRXL ( CK , D , Q , QN , RN );
    input CK ;
    input D ;
    output Q ;
    output QN ;
    input RN ;
endmodule 
module DFFX1 ( CK , D , Q , QN );
    input CK ;
    input D ;
    output Q ;
    output QN ;
endmodule 
module CLKMX2X12 ( A , B , S0 , Y );
    input A ;
    input B ;
    input S0 ;
    output Y ;
endmodule 
module CLKMX2X2 ( A , B , S0 , Y );
    input A ;
    input B ;
    input S0 ;
    output Y ;
endmodule 
module CLKMX2X3 ( A , B , S0 , Y );
    input A ;
    input B ;
    input S0 ;
    output Y ;
endmodule 
module CLKMX2X4 ( A , B , S0 , Y );
    input A ;
    input B ;
    input S0 ;
    output Y ;
endmodule 
module CLKMX2X6 ( A , B , S0 , Y );
    input A ;
    input B ;
    input S0 ;
    output Y ;
endmodule 
module CLKMX2X8 ( A , B , S0 , Y );
    input A ;
    input B ;
    input S0 ;
    output Y ;
endmodule 
module CLKXOR2X1 ( A , B , Y );
    input A ;
    input B ;
    output Y ;
endmodule 
module CLKXOR2X2 ( A , B , Y );
    input A ;
    input B ;
    output Y ;
endmodule 
module CLKXOR2X4 ( A , B , Y );
    input A ;
    input B ;
    output Y ;
endmodule 
module CLKXOR2X8 ( A , B , Y );
    input A ;
    input B ;
    output Y ;
endmodule 
module CMPR22X2 ( A , B , CO , S );
    input A ;
    input B ;
    output CO ;
    output S ;
endmodule 
module OAI2BB2X1 ( A0N , A1N , B0 , B1 , Y );
    input A0N ;
    input A1N ;
    input B0 ;
    input B1 ;
    output Y ;
endmodule 
module NOR2XL ( A , B , Y );
    input A ;
    input B ;
    output Y ;
endmodule 
module NOR3BX1 ( AN , B , C , Y );
    input AN ;
    input B ;
    input C ;
    output Y ;
endmodule 
module NOR3BX2 ( AN , B , C , Y );
    input AN ;
    input B ;
    input C ;
    output Y ;
endmodule 
module NOR3BX4 ( AN , B , C , Y );
    input AN ;
    input B ;
    input C ;
    output Y ;
endmodule 
module EDFFTRX2 ( CK , D , E , Q , QN , RN );
    input CK ;
    input D ;
    input E ;
    output Q ;
    output QN ;
    input RN ;
endmodule 
module EDFFTRX4 ( CK , D , E , Q , QN , RN );
    input CK ;
    input D ;
    input E ;
    output Q ;
    output QN ;
    input RN ;
endmodule 
module EDFFTRXL ( CK , D , E , Q , QN , RN );
    input CK ;
    input D ;
    input E ;
    output Q ;
    output QN ;
    input RN ;
endmodule 
module EDFFX1 ( CK , D , E , Q , QN );
    input CK ;
    input D ;
    input E ;
    output Q ;
    output QN ;
endmodule 
module EDFFX2 ( CK , D , E , Q , QN );
    input CK ;
    input D ;
    input E ;
    output Q ;
    output QN ;
endmodule 
module EDFFX4 ( CK , D , E , Q , QN );
    input CK ;
    input D ;
    input E ;
    output Q ;
    output QN ;
endmodule 
module EDFFXL ( CK , D , E , Q , QN );
    input CK ;
    input D ;
    input E ;
    output Q ;
    output QN ;
endmodule 
module FILL16 ();
endmodule 
module FILL1 ();
endmodule 
module FILL2 ();
endmodule 
module FILL32 ();
endmodule 
module FILL4 ();
endmodule 
module FILL64 ();
endmodule 
module DFFRHQX1 ( CK , D , Q , RN );
    input CK ;
    input D ;
    output Q ;
    input RN ;
endmodule 
module DFFRHQX2 ( CK , D , Q , RN );
    input CK ;
    input D ;
    output Q ;
    input RN ;
endmodule 
module DFFRHQX4 ( CK , D , Q , RN );
    input CK ;
    input D ;
    output Q ;
    input RN ;
endmodule 
module DFFRHQX8 ( CK , D , Q , RN );
    input CK ;
    input D ;
    output Q ;
    input RN ;
endmodule 
module DFFRX1 ( CK , D , Q , QN , RN );
    input CK ;
    input D ;
    output Q ;
    output QN ;
    input RN ;
endmodule 
module DFFRX2 ( CK , D , Q , QN , RN );
    input CK ;
    input D ;
    output Q ;
    output QN ;
    input RN ;
endmodule 
module DFFRX4 ( CK , D , Q , QN , RN );
    input CK ;
    input D ;
    output Q ;
    output QN ;
    input RN ;
endmodule 
module DFFRXL ( CK , D , Q , QN , RN );
    input CK ;
    input D ;
    output Q ;
    output QN ;
    input RN ;
endmodule 
module DFFSHQX1 ( CK , D , Q , SN );
    input CK ;
    input D ;
    output Q ;
    input SN ;
endmodule 
module DFFSHQX2 ( CK , D , Q , SN );
    input CK ;
    input D ;
    output Q ;
    input SN ;
endmodule 
module DFFSHQX4 ( CK , D , Q , SN );
    input CK ;
    input D ;
    output Q ;
    input SN ;
endmodule 
module DFFSHQX8 ( CK , D , Q , SN );
    input CK ;
    input D ;
    output Q ;
    input SN ;
endmodule 
module DFFSRHQX1 ( CK , D , Q , RN , SN );
    input CK ;
    input D ;
    output Q ;
    input RN ;
    input SN ;
endmodule 
module DFFSRHQX2 ( CK , D , Q , RN , SN );
    input CK ;
    input D ;
    output Q ;
    input RN ;
    input SN ;
endmodule 
module DFFSRHQX4 ( CK , D , Q , RN , SN );
    input CK ;
    input D ;
    output Q ;
    input RN ;
    input SN ;
endmodule 
module DFFSRHQX8 ( CK , D , Q , RN , SN );
    input CK ;
    input D ;
    output Q ;
    input RN ;
    input SN ;
endmodule 
module MX2X1 ( A , B , S0 , Y );
    input A ;
    input B ;
    input S0 ;
    output Y ;
endmodule 
module MX2X2 ( A , B , S0 , Y );
    input A ;
    input B ;
    input S0 ;
    output Y ;
endmodule 
module MX2X4 ( A , B , S0 , Y );
    input A ;
    input B ;
    input S0 ;
    output Y ;
endmodule 
module MX2X6 ( A , B , S0 , Y );
    input A ;
    input B ;
    input S0 ;
    output Y ;
endmodule 
module MX2X8 ( A , B , S0 , Y );
    input A ;
    input B ;
    input S0 ;
    output Y ;
endmodule 
module MX2XL ( A , B , S0 , Y );
    input A ;
    input B ;
    input S0 ;
    output Y ;
endmodule 
module MX3X1 ( A , B , C , S0 , S1 , Y );
    input A ;
    input B ;
    input C ;
    input S0 ;
    input S1 ;
    output Y ;
endmodule 
module MX3X2 ( A , B , C , S0 , S1 , Y );
    input A ;
    input B ;
    input C ;
    input S0 ;
    input S1 ;
    output Y ;
endmodule 
module MX3X4 ( A , B , C , S0 , S1 , Y );
    input A ;
    input B ;
    input C ;
    input S0 ;
    input S1 ;
    output Y ;
endmodule 
module MX3XL ( A , B , C , S0 , S1 , Y );
    input A ;
    input B ;
    input C ;
    input S0 ;
    input S1 ;
    output Y ;
endmodule 
module MX4X1 ( A , B , C , D , S0 , S1 , Y );
    input A ;
    input B ;
    input C ;
    input D ;
    input S0 ;
    input S1 ;
    output Y ;
endmodule 
module MX4X2 ( A , B , C , D , S0 , S1 , Y );
    input A ;
    input B ;
    input C ;
    input D ;
    input S0 ;
    input S1 ;
    output Y ;
endmodule 
module MX4X4 ( A , B , C , D , S0 , S1 , Y );
    input A ;
    input B ;
    input C ;
    input D ;
    input S0 ;
    input S1 ;
    output Y ;
endmodule 
module DFFX2 ( CK , D , Q , QN );
    input CK ;
    input D ;
    output Q ;
    output QN ;
endmodule 
module DFFX4 ( CK , D , Q , QN );
    input CK ;
    input D ;
    output Q ;
    output QN ;
endmodule 
module DFFXL ( CK , D , Q , QN );
    input CK ;
    input D ;
    output Q ;
    output QN ;
endmodule 
module DLY1X1 ( A , Y );
    input A ;
    output Y ;
endmodule 
module DLY1X4 ( A , Y );
    input A ;
    output Y ;
endmodule 
module DLY2X1 ( A , Y );
    input A ;
    output Y ;
endmodule 
module DLY2X4 ( A , Y );
    input A ;
    output Y ;
endmodule 
module DLY3X1 ( A , Y );
    input A ;
    output Y ;
endmodule 
module DLY3X4 ( A , Y );
    input A ;
    output Y ;
endmodule 
module DLY4X1 ( A , Y );
    input A ;
    output Y ;
endmodule 
module DLY4X4 ( A , Y );
    input A ;
    output Y ;
endmodule 
module EDFFHQX1 ( CK , D , E , Q );
    input CK ;
    input D ;
    input E ;
    output Q ;
endmodule 
module EDFFHQX2 ( CK , D , E , Q );
    input CK ;
    input D ;
    input E ;
    output Q ;
endmodule 
module EDFFHQX4 ( CK , D , E , Q );
    input CK ;
    input D ;
    input E ;
    output Q ;
endmodule 
module EDFFHQX8 ( CK , D , E , Q );
    input CK ;
    input D ;
    input E ;
    output Q ;
endmodule 
module EDFFTRX1 ( CK , D , E , Q , QN , RN );
    input CK ;
    input D ;
    input E ;
    output Q ;
    output QN ;
    input RN ;
endmodule 
module BUFX16 ( A , Y );
    input A ;
    output Y ;
endmodule 
module ANTENNA (A);
	input A ;
endmodule 
module AO21X1 ( A0 , A1 , B0 , Y );
    input A0 ;
    input A1 ;
    input B0 ;
    output Y ;
endmodule 
module AO21X2 ( A0 , A1 , B0 , Y );
    input A0 ;
    input A1 ;
    input B0 ;
    output Y ;
endmodule 
module AO21X4 ( A0 , A1 , B0 , Y );
    input A0 ;
    input A1 ;
    input B0 ;
    output Y ;
endmodule 
module AO21XL ( A0 , A1 , B0 , Y );
    input A0 ;
    input A1 ;
    input B0 ;
    output Y ;
endmodule 
module AO22X1 ( A0 , A1 , B0 , B1 , Y );
    input A0 ;
    input A1 ;
    input B0 ;
    input B1 ;
    output Y ;
endmodule 
module AO22X2 ( A0 , A1 , B0 , B1 , Y );
    input A0 ;
    input A1 ;
    input B0 ;
    input B1 ;
    output Y ;
endmodule 
module AO22X4 ( A0 , A1 , B0 , B1 , Y );
    input A0 ;
    input A1 ;
    input B0 ;
    input B1 ;
    output Y ;
endmodule 
module AO22XL ( A0 , A1 , B0 , B1 , Y );
    input A0 ;
    input A1 ;
    input B0 ;
    input B1 ;
    output Y ;
endmodule 
module AOI211X1 ( A0 , A1 , B0 , C0 , Y );
    input A0 ;
    input A1 ;
    input B0 ;
    input C0 ;
    output Y ;
endmodule 
module AOI211X2 ( A0 , A1 , B0 , C0 , Y );
    input A0 ;
    input A1 ;
    input B0 ;
    input C0 ;
    output Y ;
endmodule 
module AOI211X4 ( A0 , A1 , B0 , C0 , Y );
    input A0 ;
    input A1 ;
    input B0 ;
    input C0 ;
    output Y ;
endmodule 
module AOI211XL ( A0 , A1 , B0 , C0 , Y );
    input A0 ;
    input A1 ;
    input B0 ;
    input C0 ;
    output Y ;
endmodule 
module AOI21X1 ( A0 , A1 , B0 , Y );
    input A0 ;
    input A1 ;
    input B0 ;
    output Y ;
endmodule 
module AOI21X2 ( A0 , A1 , B0 , Y );
    input A0 ;
    input A1 ;
    input B0 ;
    output Y ;
endmodule 
module AOI21X4 ( A0 , A1 , B0 , Y );
    input A0 ;
    input A1 ;
    input B0 ;
    output Y ;
endmodule 
module AOI21XL ( A0 , A1 , B0 , Y );
    input A0 ;
    input A1 ;
    input B0 ;
    output Y ;
endmodule 
module INVX20 ( A , Y );
    input A ;
    output Y ;
endmodule 
module INVX2 ( A , Y );
    input A ;
    output Y ;
endmodule 
module INVX3 ( A , Y );
    input A ;
    output Y ;
endmodule 
module INVX4 ( A , Y );
    input A ;
    output Y ;
endmodule 
module INVX6 ( A , Y );
    input A ;
    output Y ;
endmodule 
module INVX8 ( A , Y );
    input A ;
    output Y ;
endmodule 
module INVXL ( A , Y );
    input A ;
    output Y ;
endmodule 
module MDFFHQX1 ( CK , D0 , D1 , Q , S0 );
    input CK ;
    input D0 ;
    input D1 ;
    output Q ;
    input S0 ;
endmodule 
module MDFFHQX2 ( CK , D0 , D1 , Q , S0 );
    input CK ;
    input D0 ;
    input D1 ;
    output Q ;
    input S0 ;
endmodule 
module MDFFHQX4 ( CK , D0 , D1 , Q , S0 );
    input CK ;
    input D0 ;
    input D1 ;
    output Q ;
    input S0 ;
endmodule 
module MDFFHQX8 ( CK , D0 , D1 , Q , S0 );
    input CK ;
    input D0 ;
    input D1 ;
    output Q ;
    input S0 ;
endmodule 
module CLKINVX8 ( A , Y );
    input A ;
    output Y ;
endmodule 
module AOI2BB1X1 ( A0N , A1N , B0 , Y );
    input A0N ;
    input A1N ;
    input B0 ;
    output Y ;
endmodule 
module AOI2BB1X2 ( A0N , A1N , B0 , Y );
    input A0N ;
    input A1N ;
    input B0 ;
    output Y ;
endmodule 
module AOI2BB1X4 ( A0N , A1N , B0 , Y );
    input A0N ;
    input A1N ;
    input B0 ;
    output Y ;
endmodule 
module AOI2BB1XL ( A0N , A1N , B0 , Y );
    input A0N ;
    input A1N ;
    input B0 ;
    output Y ;
endmodule 
module AOI2BB2X1 ( A0N , A1N , B0 , B1 , Y );
    input A0N ;
    input A1N ;
    input B0 ;
    input B1 ;
    output Y ;
endmodule 
module AOI2BB2X2 ( A0N , A1N , B0 , B1 , Y );
    input A0N ;
    input A1N ;
    input B0 ;
    input B1 ;
    output Y ;
endmodule 
module AOI2BB2X4 ( A0N , A1N , B0 , B1 , Y );
    input A0N ;
    input A1N ;
    input B0 ;
    input B1 ;
    output Y ;
endmodule 
module AOI2BB2XL ( A0N , A1N , B0 , B1 , Y );
    input A0N ;
    input A1N ;
    input B0 ;
    input B1 ;
    output Y ;
endmodule 
module AOI31X1 ( A0 , A1 , A2 , B0 , Y );
    input A0 ;
    input A1 ;
    input A2 ;
    input B0 ;
    output Y ;
endmodule 
module AOI31X2 ( A0 , A1 , A2 , B0 , Y );
    input A0 ;
    input A1 ;
    input A2 ;
    input B0 ;
    output Y ;
endmodule 
module AOI31X4 ( A0 , A1 , A2 , B0 , Y );
    input A0 ;
    input A1 ;
    input A2 ;
    input B0 ;
    output Y ;
endmodule 
module AOI31XL ( A0 , A1 , A2 , B0 , Y );
    input A0 ;
    input A1 ;
    input A2 ;
    input B0 ;
    output Y ;
endmodule 
module AOI32X1 ( A0 , A1 , A2 , B0 , B1 , Y );
    input A0 ;
    input A1 ;
    input A2 ;
    input B0 ;
    input B1 ;
    output Y ;
endmodule 
module AOI32X2 ( A0 , A1 , A2 , B0 , B1 , Y );
    input A0 ;
    input A1 ;
    input A2 ;
    input B0 ;
    input B1 ;
    output Y ;
endmodule 
module AOI32X4 ( A0 , A1 , A2 , B0 , B1 , Y );
    input A0 ;
    input A1 ;
    input A2 ;
    input B0 ;
    input B1 ;
    output Y ;
endmodule 
module AOI32XL ( A0 , A1 , A2 , B0 , B1 , Y );
    input A0 ;
    input A1 ;
    input A2 ;
    input B0 ;
    input B1 ;
    output Y ;
endmodule 
module AOI33X1 ( A0 , A1 , A2 , B0 , B1 , B2 , Y );
    input A0 ;
    input A1 ;
    input A2 ;
    input B0 ;
    input B1 ;
    input B2 ;
    output Y ;
endmodule 
module AOI33X2 ( A0 , A1 , A2 , B0 , B1 , B2 , Y );
    input A0 ;
    input A1 ;
    input A2 ;
    input B0 ;
    input B1 ;
    input B2 ;
    output Y ;
endmodule 
module AOI33X4 ( A0 , A1 , A2 , B0 , B1 , B2 , Y );
    input A0 ;
    input A1 ;
    input A2 ;
    input B0 ;
    input B1 ;
    input B2 ;
    output Y ;
endmodule 
module AOI33XL ( A0 , A1 , A2 , B0 , B1 , B2 , Y );
    input A0 ;
    input A1 ;
    input A2 ;
    input B0 ;
    input B1 ;
    input B2 ;
    output Y ;
endmodule 
module BENCX1 ( A , M0 , M1 , M2 , S , X2 );
    output A ;
    input M0 ;
    input M1 ;
    input M2 ;
    output S ;
    output X2 ;
endmodule 
module BENCX2 ( A , M0 , M1 , M2 , S , X2 );
    output A ;
    input M0 ;
    input M1 ;
    input M2 ;
    output S ;
    output X2 ;
endmodule 
module BENCX4 ( A , M0 , M1 , M2 , S , X2 );
    output A ;
    input M0 ;
    input M1 ;
    input M2 ;
    output S ;
    output X2 ;
endmodule 
module BMXIX2 ( A , M0 , M1 , PPN , S , X2 );
    input A ;
    input M0 ;
    input M1 ;
    output PPN ;
    input S ;
    input X2 ;
endmodule 
module BMXIX4 ( A , M0 , M1 , PPN , S , X2 );
    input A ;
    input M0 ;
    input M1 ;
    output PPN ;
    input S ;
    input X2 ;
endmodule 
module BMXX2 ( A , M0 , M1 , PP , S , X2 );
    input A ;
    input M0 ;
    input M1 ;
    output PP ;
    input S ;
    input X2 ;
endmodule 
module BMXX4 ( A , M0 , M1 , PP , S , X2 );
    input A ;
    input M0 ;
    input M1 ;
    output PP ;
    input S ;
    input X2 ;
endmodule 
module BUFX12 ( A , Y );
    input A ;
    output Y ;
endmodule 
module DFFQXL ( CK , D , Q );
    input CK ;
    input D ;
    output Q ;
endmodule 
module BUFX20 ( A , Y );
    input A ;
    output Y ;
endmodule 
module BUFX2 ( A , Y );
    input A ;
    output Y ;
endmodule 
module BUFX3 ( A , Y );
    input A ;
    output Y ;
endmodule 
module BUFX4 ( A , Y );
    input A ;
    output Y ;
endmodule 
module BUFX6 ( A , Y );
    input A ;
    output Y ;
endmodule 
module BUFX8 ( A , Y );
    input A ;
    output Y ;
endmodule 
module CLKAND2X12 ( A , B , Y );
    input A ;
    input B ;
    output Y ;
endmodule 
module CLKAND2X2 ( A , B , Y );
    input A ;
    input B ;
    output Y ;
endmodule 
module CLKAND2X3 ( A , B , Y );
    input A ;
    input B ;
    output Y ;
endmodule 
module CLKAND2X4 ( A , B , Y );
    input A ;
    input B ;
    output Y ;
endmodule 
module CLKAND2X6 ( A , B , Y );
    input A ;
    input B ;
    output Y ;
endmodule 
module CLKAND2X8 ( A , B , Y );
    input A ;
    input B ;
    output Y ;
endmodule 
module CLKBUFX12 ( A , Y );
    input A ;
    output Y ;
endmodule 
module CLKBUFX16 ( A , Y );
    input A ;
    output Y ;
endmodule 
module CLKBUFX20 ( A , Y );
    input A ;
    output Y ;
endmodule 
module CLKBUFX2 ( A , Y );
    input A ;
    output Y ;
endmodule 
module CLKBUFX3 ( A , Y );
    input A ;
    output Y ;
endmodule 
module CLKBUFX4 ( A , Y );
    input A ;
    output Y ;
endmodule 
module CLKBUFX6 ( A , Y );
    input A ;
    output Y ;
endmodule 
module CLKBUFX8 ( A , Y );
    input A ;
    output Y ;
endmodule 
module CLKINVX12 ( A , Y );
    input A ;
    output Y ;
endmodule 
module CLKINVX16 ( A , Y );
    input A ;
    output Y ;
endmodule 
module CLKINVX1 ( A , Y );
    input A ;
    output Y ;
endmodule 
module CLKINVX20 ( A , Y );
    input A ;
    output Y ;
endmodule 
module CLKINVX2 ( A , Y );
    input A ;
    output Y ;
endmodule 
module CLKINVX3 ( A , Y );
    input A ;
    output Y ;
endmodule 
module CLKINVX4 ( A , Y );
    input A ;
    output Y ;
endmodule 
module CLKINVX6 ( A , Y );
    input A ;
    output Y ;
endmodule 
module ADDFXL ( A , B , CI , CO , S );
    input A ;
    input B ;
    input CI ;
    output CO ;
    output S ;
endmodule 
module ADDHX1 ( A , B , CO , S );
    input A ;
    input B ;
    output CO ;
    output S ;
endmodule 
module ADDHX2 ( A , B , CO , S );
    input A ;
    input B ;
    output CO ;
    output S ;
endmodule 
module ADDHX4 ( A , B , CO , S );
    input A ;
    input B ;
    output CO ;
    output S ;
endmodule 
module ADDHXL ( A , B , CO , S );
    input A ;
    input B ;
    output CO ;
    output S ;
endmodule 
module AFCSHCINX2 ( A , B , CI0N , CI1N , CO0 , CO1 , CS , S );
    input A ;
    input B ;
    input CI0N ;
    input CI1N ;
    output CO0 ;
    output CO1 ;
    input CS ;
    output S ;
endmodule 
module AFCSHCINX4 ( A , B , CI0N , CI1N , CO0 , CO1 , CS , S );
    input A ;
    input B ;
    input CI0N ;
    input CI1N ;
    output CO0 ;
    output CO1 ;
    input CS ;
    output S ;
endmodule 
module AFCSHCONX2 ( A , B , CI0 , CI1 , CO0N , CO1N , CS , S );
    input A ;
    input B ;
    input CI0 ;
    input CI1 ;
    output CO0N ;
    output CO1N ;
    input CS ;
    output S ;
endmodule 
module AFCSHCONX4 ( A , B , CI0 , CI1 , CO0N , CO1N , CS , S );
    input A ;
    input B ;
    input CI0 ;
    input CI1 ;
    output CO0N ;
    output CO1N ;
    input CS ;
    output S ;
endmodule 
module AFCSIHCONX2 ( A , B , CO0N , CO1N , CS , S );
    input A ;
    input B ;
    output CO0N ;
    output CO1N ;
    input CS ;
    output S ;
endmodule 
module AFCSIHCONX4 ( A , B , CO0N , CO1N , CS , S );
    input A ;
    input B ;
    output CO0N ;
    output CO1N ;
    input CS ;
    output S ;
endmodule 
module AFHCINX2 ( A , B , CIN , CO , S );
    input A ;
    input B ;
    input CIN ;
    output CO ;
    output S ;
endmodule 
module CMPR22X4 ( A , B , CO , S );
    input A ;
    input B ;
    output CO ;
    output S ;
endmodule 
module CMPR32X2 ( A , B , C , CO , S );
    input A ;
    input B ;
    input C ;
    output CO ;
    output S ;
endmodule 
module CMPR32X4 ( A , B , C , CO , S );
    input A ;
    input B ;
    input C ;
    output CO ;
    output S ;
endmodule 
module CMPR42X1 ( A , B , C , CO , D , ICI , ICO , S );
    input A ;
    input B ;
    input C ;
    output CO ;
    input D ;
    input ICI ;
    output ICO ;
    output S ;
endmodule 
module CMPR42X2 ( A , B , C , CO , D , ICI , ICO , S );
    input A ;
    input B ;
    input C ;
    output CO ;
    input D ;
    input ICI ;
    output ICO ;
    output S ;
endmodule 
module CMPR42X4 ( A , B , C , CO , D , ICI , ICO , S );
    input A ;
    input B ;
    input C ;
    output CO ;
    input D ;
    input ICI ;
    output ICO ;
    output S ;
endmodule 
module DFFHQX1 ( CK , D , Q );
    input CK ;
    input D ;
    output Q ;
endmodule 
module DFFHQX2 ( CK , D , Q );
    input CK ;
    input D ;
    output Q ;
endmodule 
module DFFHQX4 ( CK , D , Q );
    input CK ;
    input D ;
    output Q ;
endmodule 
module DFFHQX8 ( CK , D , Q );
    input CK ;
    input D ;
    output Q ;
endmodule 
module DFFNSRX1 ( CKN , D , Q , QN , RN , SN );
    input CKN ;
    input D ;
    output Q ;
    output QN ;
    input RN ;
    input SN ;
endmodule 
module DFFNSRX2 ( CKN , D , Q , QN , RN , SN );
    input CKN ;
    input D ;
    output Q ;
    output QN ;
    input RN ;
    input SN ;
endmodule 
module DFFNSRX4 ( CKN , D , Q , QN , RN , SN );
    input CKN ;
    input D ;
    output Q ;
    output QN ;
    input RN ;
    input SN ;
endmodule 
module DFFNSRXL ( CKN , D , Q , QN , RN , SN );
    input CKN ;
    input D ;
    output Q ;
    output QN ;
    input RN ;
    input SN ;
endmodule 
module DFFQX1 ( CK , D , Q );
    input CK ;
    input D ;
    output Q ;
endmodule 
module DFFQX2 ( CK , D , Q );
    input CK ;
    input D ;
    output Q ;
endmodule 
module DFFQX4 ( CK , D , Q );
    input CK ;
    input D ;
    output Q ;
endmodule 
module AND3X1 ( A , B , C , Y );
    input A ;
    input B ;
    input C ;
    output Y ;
endmodule 
module AND3X2 ( A , B , C , Y );
    input A ;
    input B ;
    input C ;
    output Y ;
endmodule 
module AND3X4 ( A , B , C , Y );
    input A ;
    input B ;
    input C ;
    output Y ;
endmodule 
module AND3X6 ( A , B , C , Y );
    input A ;
    input B ;
    input C ;
    output Y ;
endmodule 
module AND3X8 ( A , B , C , Y );
    input A ;
    input B ;
    input C ;
    output Y ;
endmodule 
module AND3XL ( A , B , C , Y );
    input A ;
    input B ;
    input C ;
    output Y ;
endmodule 
module AND4X1 ( A , B , C , D , Y );
    input A ;
    input B ;
    input C ;
    input D ;
    output Y ;
endmodule 
module AND4X2 ( A , B , C , D , Y );
    input A ;
    input B ;
    input C ;
    input D ;
    output Y ;
endmodule 
module AND4X4 ( A , B , C , D , Y );
    input A ;
    input B ;
    input C ;
    input D ;
    output Y ;
endmodule 
module AND4X6 ( A , B , C , D , Y );
    input A ;
    input B ;
    input C ;
    input D ;
    output Y ;
endmodule 
module AND4X8 ( A , B , C , D , Y );
    input A ;
    input B ;
    input C ;
    input D ;
    output Y ;
endmodule 
module AND4XL ( A , B , C , D , Y );
    input A ;
    input B ;
    input C ;
    input D ;
    output Y ;
endmodule 
module ACCSHCINX2 ( A , B , CI0N , CI1N , CO0 , CO1 );
    input A ;
    input B ;
    input CI0N ;
    input CI1N ;
    output CO0 ;
    output CO1 ;
endmodule 
module ACCSHCINX4 ( A , B , CI0N , CI1N , CO0 , CO1 );
    input A ;
    input B ;
    input CI0N ;
    input CI1N ;
    output CO0 ;
    output CO1 ;
endmodule 
module ACCSHCONX2 ( A , B , CI0 , CI1 , CO0N , CO1N );
    input A ;
    input B ;
    input CI0 ;
    input CI1 ;
    output CO0N ;
    output CO1N ;
endmodule 
module ACCSHCONX4 ( A , B , CI0 , CI1 , CO0N , CO1N );
    input A ;
    input B ;
    input CI0 ;
    input CI1 ;
    output CO0N ;
    output CO1N ;
endmodule 
module ACCSIHCONX2 ( A , B , CO0N , CO1N );
    input A ;
    input B ;
    output CO0N ;
    output CO1N ;
endmodule 
module ACCSIHCONX4 ( A , B , CO0N , CO1N );
    input A ;
    input B ;
    output CO0N ;
    output CO1N ;
endmodule 
module ACHCINX2 ( A , B , CIN , CO );
    input A ;
    input B ;
    input CIN ;
    output CO ;
endmodule 
module ACHCINX4 ( A , B , CIN , CO );
    input A ;
    input B ;
    input CIN ;
    output CO ;
endmodule 
module ACHCONX2 ( A , B , CI , CON );
    input A ;
    input B ;
    input CI ;
    output CON ;
endmodule 
module ACHCONX4 ( A , B , CI , CON );
    input A ;
    input B ;
    input CI ;
    output CON ;
endmodule 
module ADDFHX1 ( A , B , CI , CO , S );
    input A ;
    input B ;
    input CI ;
    output CO ;
    output S ;
endmodule 
module ADDFHX2 ( A , B , CI , CO , S );
    input A ;
    input B ;
    input CI ;
    output CO ;
    output S ;
endmodule 
module ADDFHX4 ( A , B , CI , CO , S );
    input A ;
    input B ;
    input CI ;
    output CO ;
    output S ;
endmodule 
module ADDFHXL ( A , B , CI , CO , S );
    input A ;
    input B ;
    input CI ;
    output CO ;
    output S ;
endmodule 
module ADDFX1 ( A , B , CI , CO , S );
    input A ;
    input B ;
    input CI ;
    output CO ;
    output S ;
endmodule 
module ADDFX2 ( A , B , CI , CO , S );
    input A ;
    input B ;
    input CI ;
    output CO ;
    output S ;
endmodule 
module ADDFX4 ( A , B , CI , CO , S );
    input A ;
    input B ;
    input CI ;
    output CO ;
    output S ;
endmodule 
module AOI221X1 ( A0 , A1 , B0 , B1 , C0 , Y );
    input A0 ;
    input A1 ;
    input B0 ;
    input B1 ;
    input C0 ;
    output Y ;
endmodule 
module AOI221X2 ( A0 , A1 , B0 , B1 , C0 , Y );
    input A0 ;
    input A1 ;
    input B0 ;
    input B1 ;
    input C0 ;
    output Y ;
endmodule 
module AOI221X4 ( A0 , A1 , B0 , B1 , C0 , Y );
    input A0 ;
    input A1 ;
    input B0 ;
    input B1 ;
    input C0 ;
    output Y ;
endmodule 
module AOI221XL ( A0 , A1 , B0 , B1 , C0 , Y );
    input A0 ;
    input A1 ;
    input B0 ;
    input B1 ;
    input C0 ;
    output Y ;
endmodule 
module AOI222X1 ( A0 , A1 , B0 , B1 , C0 , C1 , Y );
    input A0 ;
    input A1 ;
    input B0 ;
    input B1 ;
    input C0 ;
    input C1 ;
    output Y ;
endmodule 
module AOI222X2 ( A0 , A1 , B0 , B1 , C0 , C1 , Y );
    input A0 ;
    input A1 ;
    input B0 ;
    input B1 ;
    input C0 ;
    input C1 ;
    output Y ;
endmodule 
module AOI222X4 ( A0 , A1 , B0 , B1 , C0 , C1 , Y );
    input A0 ;
    input A1 ;
    input B0 ;
    input B1 ;
    input C0 ;
    input C1 ;
    output Y ;
endmodule 
module AOI222XL ( A0 , A1 , B0 , B1 , C0 , C1 , Y );
    input A0 ;
    input A1 ;
    input B0 ;
    input B1 ;
    input C0 ;
    input C1 ;
    output Y ;
endmodule 
module AOI22X1 ( A0 , A1 , B0 , B1 , Y );
    input A0 ;
    input A1 ;
    input B0 ;
    input B1 ;
    output Y ;
endmodule 
module AOI22X2 ( A0 , A1 , B0 , B1 , Y );
    input A0 ;
    input A1 ;
    input B0 ;
    input B1 ;
    output Y ;
endmodule 
module AOI22X4 ( A0 , A1 , B0 , B1 , Y );
    input A0 ;
    input A1 ;
    input B0 ;
    input B1 ;
    output Y ;
endmodule 
module AOI22XL ( A0 , A1 , B0 , B1 , Y );
    input A0 ;
    input A1 ;
    input B0 ;
    input B1 ;
    output Y ;
endmodule 
module AFHCINX4 ( A , B , CIN , CO , S );
    input A ;
    input B ;
    input CIN ;
    output CO ;
    output S ;
endmodule 
module AFHCONX2 ( A , B , CI , CON , S );
    input A ;
    input B ;
    input CI ;
    output CON ;
    output S ;
endmodule 
module AFHCONX4 ( A , B , CI , CON , S );
    input A ;
    input B ;
    input CI ;
    output CON ;
    output S ;
endmodule 
module AHCSHCINX2 ( A , CIN , CO , CS , S );
    input A ;
    input CIN ;
    output CO ;
    input CS ;
    output S ;
endmodule 
module AHCSHCINX4 ( A , CIN , CO , CS , S );
    input A ;
    input CIN ;
    output CO ;
    input CS ;
    output S ;
endmodule 
module AHCSHCONX2 ( A , CI , CON , CS , S );
    input A ;
    input CI ;
    output CON ;
    input CS ;
    output S ;
endmodule 
module AHCSHCONX4 ( A , CI , CON , CS , S );
    input A ;
    input CI ;
    output CON ;
    input CS ;
    output S ;
endmodule 
module AHHCINX2 ( A , CIN , CO , S );
    input A ;
    input CIN ;
    output CO ;
    output S ;
endmodule 
module AHHCINX4 ( A , CIN , CO , S );
    input A ;
    input CIN ;
    output CO ;
    output S ;
endmodule 
module AHHCONX2 ( A , CI , CON , S );
    input A ;
    input CI ;
    output CON ;
    output S ;
endmodule 
module AHHCONX4 ( A , CI , CON , S );
    input A ;
    input CI ;
    output CON ;
    output S ;
endmodule 
module AND2X1 ( A , B , Y );
    input A ;
    input B ;
    output Y ;
endmodule 
module AND2X2 ( A , B , Y );
    input A ;
    input B ;
    output Y ;
endmodule 
module AND2X4 ( A , B , Y );
    input A ;
    input B ;
    output Y ;
endmodule 
module AND2X6 ( A , B , Y );
    input A ;
    input B ;
    output Y ;
endmodule 
module AND2X8 ( A , B , Y );
    input A ;
    input B ;
    output Y ;
endmodule 
module AND2XL ( A , B , Y );
    input A ;
    input B ;
    output Y ;
endmodule 

