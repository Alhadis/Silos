module XOR2X1 (IN1,IN2,Q);
	input IN1,IN2
	output Q
endmodule


module AND2X1 (IN1,IN2,Q);
	input IN1,IN2
	output Q
endmodule


module AO22X1 (IN1,IN2,IN3,IN4,Q);
	input IN1,IN2,IN3,IN4
	output Q
endmodule



module OAI21X1 (IN1,IN2,IN3,QN);
	input IN1,IN2,IN3
	output QN
endmodule



module AOI21X1 (IN1,IN2,IN3,QN);
	input IN1,IN2,IN3
	output QN
endmodule


module OR3X1 (IN1,IN2,IN3,Q);
	input IN1,IN2,IN3
	output Q
endmodule



module OR2X1 (IN1,IN2,Q);
	input IN1,IN2
	output Q
endmodule


module OA221X1 (IN1,IN2,IN3,IN4,IN5,Q);
	input IN1,IN2,IN3,IN4,IN5
	output Q
endmodule



module NOR3X0 (IN1,IN2,IN3,QN);
	input IN1,IN2,IN3
	output QN
endmodule



module AOI22X1 (IN1,IN2,IN3,IN4,QN);
	input IN1,IN2,IN3,IN4
	output QN
endmodule





module OA22X1 (IN1,IN2,IN3,IN4,Q);
	input IN1,IN2,IN3,IN4
	output Q
endmodule




module NOR2X0 (IN1,IN2,QN);
	input IN1,IN2
	output QN
endmodule


module OA21X1 (IN1,IN2,IN3,Q);
	input IN1,IN2,IN3
	output Q
endmodule




module AND3X1 (IN1,IN2,IN3,Q);
	input IN1,IN2,IN3
	output Q
endmodule



module NAND3X0 (IN1,IN2,IN3,QN);
	input IN1,IN2,IN3
	output QN
endmodule


module XNOR2X1 (IN1,IN2,Q);
	input IN1,IN2
	output Q
endmodule



module INVX0 (INP,ZN);
	input INP
	output ZN
endmodule



module OAI22X1 (IN1,IN2,IN3,IN4,QN);
	input IN1,IN2,IN3,IN4
	output QN
endmodule



module NAND2X0 (IN1,IN2,QN);
	input IN1,IN2
	output QN
endmodule








































