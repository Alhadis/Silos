`timescale 1ns/1ps
`include "pckg_block.vh"
// Блок коммутации и формирования пакета для передачи на LVDS канал
module pckg_block(
    input wire clk,
    // Запуск устройства
    input wire start,

    // Порты чтения из FIFO
    output wire rd_en_fifo_1,
    input wire [`BUFF_SIZE-1:0] dat_from_fifo_1,
    output wire rd_en_fifo_2,
    input wire [`BUFF_SIZE-1:0] dat_from_fifo_2,
    // Связь с блоком управления
    // Готовность принимать следующий пакет
    output wire next,
    // Выбор приёмного канала. Кодировка:
    input wire [1:0] rdy_cnl,              // 0 - Передаем пустой пакет
    // 1 - Передаём данный из fifo_1
    // 2 - Передаём данные из fifo_2
    // Интерфейс передатчика LVDS
    // Флаг, сообщающий, что передатчик занят
    input wire tx_busy,
    // Данные для передачи
    output wire [`CH_NUM*`BUFF_SIZE-1:0] data_out,
    // Флаг готовности данных для передачи
    output wire tx_ena
);
    parameter st_start = 4'b0000, st_h1 = 4'b0001, st_empty_pck = 4'b0010, st_size = 4'b0011, st_tx_fifo_1 = 4'b0100, st_tx_fifo_2 = 4'b0101, st_tail = 4'b0110, st_next = 4'b1000; //Объявляем и кодируем автомат состояний для приёмника
    parameter size_data = `DATA_BYTES_SIZE; // Количество байт данных
    parameter size_signals = `BUFF_SIZE-1; 	// Разрядность источников сигнала
    parameter [7:0] tail = 8'h8F;			// байт-конец сообщения
	reg [4:0] st = st_start;    // Начальное состояние
    // Объявляем сигналы
    reg rd_en_1 = 1'b0;
    reg rd_en_2 = 1'b0;
    reg next_i = 1'b0;
    // Счётчик колличества слов в пакете
    reg [3:0] cnt_size = 4'h0;
    // Счётчик для сборки целого байта
    reg [2:0] cnt_byte = 3'b000;
    // СИгналы для вывода наружу
    reg tx_ena_i = 1'b0;
    reg [`CH_NUM*`BUFF_SIZE-1:0] data_out_i = 8'b0;
    // Вывод наружу
    assign data_out = data_out_i;
    assign next = next_i;

    assign rd_en_fifo_1 = rd_en_1;
    assign rd_en_fifo_2 = rd_en_2;
    
    assign tx_ena = tx_ena_i;

    // Процесс в виде цифрового автомата в котором формируется пакет,  коммутируется входной канал и отправляет данные на отправку.
    always @(posedge clk)
        begin
            case (st)
                //////////////////////////////////////////////////////////////////////////////////////////////////////////////////
                // начальное состояние. Ждём запуска устройства
                //////////////////////////////////////////////////////////////////////////////////////////////////////////////////
                st_start:
                    if (start)
                        st <= st_h1;
                //////////////////////////////////////////////////////////////////////////////////////////////////////////////////
                // Состояние передачи первого байта заголовка
                //////////////////////////////////////////////////////////////////////////////////////////////////////////////////
                st_h1:
                    // Если передатчик свободен, то отправляем на него FN, Где N - номер канала равный 2.
                    begin
                        if (tx_busy == 0)
                            begin
                                tx_ena_i <= 1;
                                data_out_i <= `HEADER_VALUE;
                                // Если код канала 0, то переходим в состояние передачи нулевого размера для пустого пакета
                                if (rdy_cnl == 0)
                                    st <= st_empty_pck;
                                    // Иначе переходим в состояние передачи размера пакета данных равным size_data байт
                                else
                                    st <= st_size;
                            end
                        else
                            tx_ena_i <= 0;
                        next_i <= 0;
                    end

                //////////////////////////////////////////////////////////////////////////////////////////////////////////////////
                // Состояние предачи нулевого размера при пустом пакете
                //////////////////////////////////////////////////////////////////////////////////////////////////////////////////
                st_empty_pck:
                    if (tx_busy == 0)
                        begin
                            tx_ena_i <= 1;
                            data_out_i <= 24'h00;
                            st <= st_next;
                        end
                    else
                        tx_ena_i <= 0;
                //////////////////////////////////////////////////////////////////////////////////////////////////////////////////
                // Передаём размер данных size_data = `DATA_BYTES_SIZE
                //////////////////////////////////////////////////////////////////////////////////////////////////////////////////
                st_size:
                    if (tx_busy == 1'b0)
                        begin
                            tx_ena_i <= 1'b1;
                            data_out_i <= size_data;
                            // Формируем пакет с даннными из фифо 1
                            if (rdy_cnl == 1)
                                st <= st_tx_fifo_1; // Следующее состояние
                                // Формируем пакет с даннми из фифо 2
                            else if (rdy_cnl == 2)
                                st <= st_tx_fifo_2; // Следующее состояние
                        end
                    else
                        tx_ena_i <= 0;

                //////////////////////////////////////////////////////////////////////////////////////////////////////////////////
                // Состояние передачи пакета данных из fifo_1 (4)
                //////////////////////////////////////////////////////////////////////////////////////////////////////////////////
                st_tx_fifo_1:
                    `send_message(dat_from_fifo_1,rd_en_1)

                //////////////////////////////////////////////////////////////////////////////////////////////////////////////////
                // Состояние передачи пакета данных из fifo_2 (5)
                //////////////////////////////////////////////////////////////////////////////////////////////////////////////////
                st_tx_fifo_2:
                    `send_message(dat_from_fifo_2,rd_en_2)
				st_tail:
					if (tx_busy == 0)
                        begin
                            tx_ena_i <= 1;
                            data_out_i <= tail;
                            st <= st_next;
                        end
                    else
                        tx_ena_i <= 0;
                
				//////////////////////////////////////////////////////////////////////////////////////////////////////////////////
                // Состояние конца передачи пакета. ЗАпрашиваем данне для следующего пакета.
                //////////////////////////////////////////////////////////////////////////////////////////////////////////////////
                st_next:
                    begin
					if (tx_busy == 0)
						tx_ena_i <= 1;
                    else
						begin
                        tx_ena_i <= 0;
                        next_i <= 1;
                        st <= st_h1;
						end
                    end

            endcase
        end
endmodule: pckg_block