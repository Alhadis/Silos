module winreg

// TODO Implement.