

module Store(CLOCK_50);
//***************************************************************
input CLOCK_50;
reg [31:0] dataMemory; // data memory buffer
//***************************************************************

/* recieve result and address */
/* access data memory pointer to send information information */


endmodule