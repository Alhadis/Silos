module design(I1,I2,I3,I4,I5,I6,I7,I8,I9,I10,I11,I12,I13,I14,I15,I16,I17,I18,I19,I20,
I21,I22,I23,I24,I25,I26,I27,I28,I29,I30,I31,I32,I33,I34,I35,I36,I37,I38,I39,I40,I41,
I42,I43,I44,I45,I46,I47,I48,I49,I50,I51,I52,I53,I54,I55,I56,I57,I58,I59,I60,I61,I62,
I63,I64,I65,I66,I67,I68,I69,I70,I71,I72,I73,I74,I75,I76,I77,I78,I79,I80,I81,I82,I83,
I84,I85,I86,I87,I88,I89,I90,I91,I92,I93,I94,I95,I96,I97,I98,I99,I100,I101,I102,I103,I104,
I105,I106,I107,I108,I109,I110,I111,I112,I113,I114,I115,I116,I117,I118,I119,I120,I121,I122,I123,I124,I125,
I126,I127,I128,I129,I130,I131,I132,I133,I134,I135,I136,I137,I138,I139,I140,I141,I142,I143,I144,I145,I146,
I147,I148,I149,I150,I151,I152,I153,I154,I155,I156,I157,I158,I159,I160,I161,I162,I163,I164,I165,I166,I167,
I168,I169,I170,I171,I172,I173,I174,I175,I176,I177,I178,I179,I180,I181,I182,I183,I184,I185,I186,I187,I188,
I189,I190,I191,I192,I193,I194,I195,I196,I197,I198,I199,I200,I201,I202,I203,I204,I205,I206,I207,I208,I209,
I210,I211,I212,I213,I214,I215,I216,I217,I218,I219,I220,I221,I222,I223,I224,I225,I226,I227,I228,I229,I230,
I231,I232,I233,I234,I235,I236,I237,I238,I239,I240,I241,I242,I243,I244,I245,I246,I247,I248,I249,I250,I251,
I252,I253,I254,I255,I256,I257,I258,I259,I260,I261,I262,I263,I264,I265,I266,I267,I268,I269,I270,I271,I272,
I273,I274,I275,I276,I277,I278,I279,I280,I281,I282,I283,I284,I285,I286,I287,I288,I289,I290,I291,I292,I293,
I294,I295,I296,I297,I298,I299,I300,I301,I302,I303,I304,I305,I306,I307,I308,I309,I310,I311,I312,I313,I314,
I315,I316,I317,I318,I319,I320,I321,I322,I323,I324,I325,I326,I327,I328,I329,I330,I331,I332,I333,I334,I335,
I336,I337,I338,I339,I340,I341,I342,I343,I344,I345,I346,I347,I348,I349,I350,I351,I352,I353,I354,I355,I356,
I357,I358,I359,I360,I361,I362,I363,I364,I365,I366,I367,I368,I369,I370,I371,I372,I373,I374,I375,I376,I377,
I378,I379,I380,I381,I382,I383,I384,I385,I386,I387,I388,I389,I390,I391,I392,I393,I394,I395,I396,I397,I398,
I399,I400,I401,I402,I403,I404,I405,I406,I407,I408,I409,I410,I411,I412,I413,I414,I415,I416,I417,I418,I419,
I420,I421,I422,I423,I424,I425,I426,I427,I428,I429,I430,I431,I432,I433,I434,I435,I436,I437,I438,I439,I440,
I441,I442,I443,I444,I445,I446,I447,I448,I449,I450,I451,I452,I453,I454,I455,I456,I457,I458,I459,I460,I461,
I462,I463,I464,I465,I466,I467,I468,I469,I470,I471,I472,I473,I474,I475,I476,I477,I478,I479,I480,I481,I482,
I483,I484,I485,I486,I487,I488,I489,I490,I491,I492,I493,I494,I495,I496,I497,I498,I499,I500,I501,I502,I503,
I504,I505,I506,I507,I508,I509,I510,I511,I512,I513,I514,I515,I516,I517,I518,I519,I520,I521,I522,I523,I524,
I525,I526,I527,I528,I529,I530,I531,I532,I533,I534,I535,I536,I537,I538,I539,I540,I541,I542,I543,I544,I545,
I546,I547,I548,I549,I550,I551,I552,I553,I554,I555,I556,I557,I558,I559,I560,I561,I562,I563,I564,I565,I566,
I567,I568,I569,I570,I571,I572,I573,I574,I575,I576,I577,I578,I579,I580,I581,I582,I583,I584,I585,I586,I587,
I588,I589,I590,I591,I592,I593,I594,I595,I596,I597,I598,I599,I600,I601,I602,I603,I604,I605,I606,I607,I608,
I609,I610,I611,I612,I613,I614,I615,I616,I617,I618,I619,I620,I621,I622,I623,I624,I625,I626,I627,I628,I629,
I630,I631,I632,I633,I634,I635,I636,I637,I638,I639,I640,I641,I642,I643,I644,I645,I646,I647,I648,I649,I650,
I651,I652,I653,I654,I655,I656,I657,I658,I659,I660,I661,I662,I663,I664,I665,I666,I667,I668,I669,I670,I671,
I672,I673,I674,I675,I676,I677,I678,I679,I680,I681,I682,I683,I684,I685,I686,I687,I688,I689,I690,I691,I692,
I693,I694,I695,I696,I697,I698,I699,I700,I701,I702,I703,I704,I705,I706,I707,I708,I709,I710,I711,I712,I713,
I714,I715,I716,I717,I718,I719,I720,I721,I722,I723,I724,I725,I726,I727,I728,I729,I730,I731,I732,I733,I734,
I735,I736,I737,I738,I739,I740,I741,I742,I743,I744,I745,I746,I747,I748,I749,I750,I751,I752,I753,I754,I755,
I756,I757,I758,I759,I760,I761,I762,I763,I764,I765,I766,I767,I768,I769,I770,I771,I772,I773,I774,I775,I776,
I777,I778,I779,I780,I781,I782,I783,I784,I785,I786,I787,I788,I789,I790,I791,I792,I793,I794,I795,I796,I797,
I798,I799,I800,I801,I802,I803,I804,I805,I806,I807,I808,I809,I810,I811,I812,I813,I814,I815,I816,I817,I818,
I819,I820,I821,I822,I823,I824,I825,I826,I827,I828,I829,I830,I831,I832,I833,I834,I835,I836,I837,I838,I839,
I840,I841,I842,I843,I844,I845,I846,I847,I848,I849,I850,I851,I852,I853,I854,I855,I856,I857,I858,I859,I860,
I861,I862,I863,I864,I865,I866,I867,I868,I869,I870,I871,I872,I873,I874,I875,I876,I877,I878,I879,I880,I881,
I882,I883,I884,I885,I886,I887,I888,I889,I890,I891,I892,I893,I894,I895,I896,I897,I898,I899,I900,I901,I902,
I903,I904,I905,I906,I907,I908,I909,I910,I911,I912,I913,I914,I915,I916,I917,I918,I919,I920,I921,I922,I923,
I924,I925,I926,I927,I928,I929,I930,I931,I932,I933,I934,I935,I936,I937,I938,I939,I940,I941,I942,I943,I944,
I945,I946,I947,I948,I949,I950,I951,I952,I953,I954,I955,I956,I957,I958,I959,I960,I961,I962,I963,I964,I965,
I966,I967,I968,I969,I970,I971,I972,I973,I974,I975,I976,I977,I978,I979,I980,I981,I982,I983,I984,I985,I986,
I987,I988,I989,I990,I991,I992,I993,I994,I995,I996,I997,I998,I999,I1000,I1001,I1002,I1003,I1004,I1005,I1006,I1007,
I1008,I1009,I1010,I1011,I1012,I1013,I1014,I1015,I1016,I1017,I1018,I1019,I1020,I1021,I1022,I1023,I1024,I1025,I1026,I1027,I1028,
I1029,I1030,I1031,I1032,I1033,I1034,I1035,I1036,I1037,I1038,I1039,I1040,I1041,I1042,I1043,I1044,I1045,I1046,I1047,I1048,I1049,
I1050,I1051,I1052,I1053,I1054,I1055,I1056,I1057,I1058,I1059,I1060,I1061,I1062,I1063,I1064,I1065,I1066,I1067,I1068,I1069,I1070,
I1071,I1072,I1073,I1074,I1075,I1076,I1077,I1078,I1079,I1080,I1081,I1082,I1083,I1084,I1085,I1086,I1087,I1088,I1089,I1090,I1091,
I1092,I1093,I1094,I1095,I1096,I1097,I1098,I1099,I1100,I1101,I1102,I1103,I1104,I1105,I1106,I1107,I1108,I1109,I1110,I1111,I1112,
I1113,I1114,I1115,I1116,I1117,I1118,I1119,I1120,I1121,I1122,I1123,I1124,I1125,I1126,I1127,I1128,I1129,I1130,I1131,I1132,I1133,
I1134,I1135,I1136,I1137,I1138,I1139,I1140,I1141,I1142,I1143,I1144,I1145,I1146,I1147,I1148,I1149,I1150,I1151,I1152,I1153,I1154,
I1155,I1156,I1157,I1158,I1159,I1160,I1161,I1162,I1163,I1164,I1165,I1166,I1167,I1168,I1169,I1170,I1171,I1172,I1173,I1174,I1175,
I1176,I1177,I1178,I1179,I1180,I1181,I1182,I1183,I1184,I1185,I1186,I1187,I1188,I1189,I1190,I1191,I1192,I1193,I1194,I1195,I1196,
I1197,I1198,I1199,I1200,I1201,I1202,I1203,I1204,I1205,I1206,I1207,I1208,I1209,I1210,I1211,I1212,I1213,I1214,I1215,I1216,I1217,
I1218,I1219,I1220,I1221,I1222,I1223,I1224,I1225,I1226,I1227,I1228,I1229,I1230,I1231,I1232,I1233,I1234,I1235,I1236,I1237,I1238,
I1239,I1240,I1241,I1242,I1243,I1244,I1245,I1246,I1247,I1248,I1249,I1250,I1251,I1252,I1253,I1254,I1255,I1256,I1257,I1258,I1259,
I1260,I1261,I1262,I1263,I1264,I1265,I1266,I1267,I1268,I1269,I1270,I1271,I1272,I1273,I1274,I1275,I1276,I1277,I1278,I1279,I1280,
I1281,I1282,I1283,I1284,I1285,I1286,I1287,I1288,I1289,I1290,I1291,I1292,I1293,I1294,I1295,I1296,I1297,I1298,I1299,I1300,I1301,
I1302,I1303,I1304,I1305,I1306,I1307,I1308,I1309,I1310,I1311,I1312,I1313,I1314,I1315,I1316,I1317,I1318,I1319,I1320,I1321,I1322,
I1323,I1324,I1325,I1326,I1327,I1328,I1329,I1330,I1331,I1332,I1333,I1334,I1335,I1336,I1337,I1338,I1339,I1340,I1341,I1342,I1343,
I1344,I1345,I1346,I1347,I1348,I1349,I1350,I1351,I1352,I1353,I1354,I1355,I1356,I1357,I1358,I1359,I1360,I1361,I1362,I1363,I1364,
I1365,I1366,I1367,I1368,I1369,I1370,I1371,I1372,I1373,I1374,I1375,I1376,I1377,I1378,I1379,I1380,I1381,I1382,I1383,I1384,I1385,
I1386,I1387,I1388,I1389,I1390,I1391,I1392,I1393,I1394,I1395,I1396,I1397,I1398,I1399,I1400,I1401,I1402,I1403,I1404,I1405,I1406,
I1407,I1408,I1409,I1410,I1411,I1412,I1413,I1414,I1415,I1416,I1417,I1418,I1419,I1420,I1421,I1422,I1423,I1424,I1425,I1426,I1427,
I1428,I1429,I1430,I1431,I1432,I1433,I1434,I1435,I1436,I1437,I1438,I1439,I1440,I1441,I1442,I1443,I1444,I1445,I1446,I1447,I1448,
I1449,I1450,I1451,I1452,I1453,I1454,I1455,I1456,I1457,I1458,I1459,I1460,I1461,I1462,I1463,I1464,I1465,I1466,I1467,I1468,I1469,
I1470,I1471,I1472,I1473,I1474,I1475,I1476,I1477,I1478,I1479,I1480,I1481,I1482,I1483,I1484,I1485,I1486,I1487,I1488,I1489,I1490,
I1491,I1492,I1493,I1494,I1495,I1496,I1497,I1498,I1499,I1500,I1501,I1502,I1503,I1504,I1505,I1506,I1507,I1508,I1509,I1510,I1511,
I1512,I1513,I1514,I1515,I1516,I1517,I1518,I1519,I1520,I1521,I1522,I1523,I1524,I1525,I1526,I1527,I1528,I1529,I1530,I1531,I1532,
I1533,I1534,I1535,I1536,I1537,I1538,I1539,I1540,I1541,I1542,I1543,I1544,I1545,I1546,I1547,I1548,I1549,I1550,I1551,I1552,I1553,
I1554,I1555,I1556,I1557,I1558,I1559,I1560,I1561,I1562,I1563,I1564,I1565,I1566,I1567,I1568,I1569,I1570,I1571,I1572,I1573,I1574,
I1575,I1576,I1577,I1578,I1579,I1580,I1581,I1582,I1583,I1584,I1585,I1586,I1587,I1588,I1589,I1590,I1591,I1592,I1593,I1594,I1595,
I1596,I1597,I1598,I1599,I1600,I1601,I1602,I1603,I1604,I1605,I1606,I1607,I1608,I1609,I1610,I1611,I1612,I1613,I1614,I1615,I1616,
I1617,I1618,I1619,I1620,I1621,I1622,I1623,I1624,I1625,I1626,I1627,I1628,I1629,I1630,I1631,I1632,I1633,I1634,I1635,I1636,I1637,
I1638,I1639,I1640,I1641,I1642,I1643,I1644,O1,O2,O3,O4,O5,O6,O7,O8,O9,O10,O11,O12,O13,O14,O15,O16,O17,O18,O19,O20,
O21,O22,O23,O24,O25,O26,O27,O28,O29,O30,O31,O32,O33,O34,O35,O36,O37,O38,O39,O40,O41,
O42,O43,O44,O45,O46,O47,O48,O49,O50,O51,O52,O53,O54,O55,O56,O57,O58,O59,O60,O61,O62,
O63,O64,O65,O66,O67,O68,O69,O70,O71,O72,O73,O74,O75,O76,O77,O78,O79,O80,O81,O82,O83,
O84,O85,O86,O87,O88,O89,O90,O91,O92,O93,O94,O95,O96,O97,O98,O99,O100,O101,O102,O103,O104,
O105,O106,O107,O108,O109,O110,O111,O112,O113,O114,O115,O116,O117,O118,O119,O120,O121,O122,O123,O124,O125,
O126,O127,O128,O129,O130,O131,O132,O133,O134,O135,O136,O137,O138,O139,O140,O141,O142,O143,O144,O145,O146,
O147,O148,O149,O150,O151,O152,O153,O154,O155,O156,O157,O158,O159,O160,O161,O162,O163,O164,O165,O166,O167,
O168,O169,O170,O171,O172,O173,O174,O175,O176,O177,O178,O179,O180,O181,O182,O183,O184,O185,O186,O187,O188,
O189,O190,O191,O192,O193,O194,O195,O196,O197,O198,O199,O200,O201,O202,O203,O204,O205,O206,O207,O208,O209,
O210,O211,O212,O213,O214,O215,O216,O217,O218,O219,O220,O221,O222,O223,O224,O225,O226,O227,O228,O229,O230,
O231,O232,O233,O234,O235,O236,O237,O238,O239,O240,O241,O242,O243,O244,O245,O246,O247,O248,O249,O250,O251,
O252,O253,O254,O255,O256,O257,O258,O259,O260,O261,O262,O263,O264,O265,O266,O267,O268,O269,O270,O271,O272,
O273,O274,O275,O276,O277,O278,O279,O280,O281,O282,O283,O284,O285,O286,O287,O288,O289,O290,O291,O292,O293,
O294,O295,O296,O297,O298,O299,O300,O301,O302,O303,O304,O305,O306,O307,O308,O309,O310,O311,O312,O313,O314,
O315,O316,O317,O318,O319,O320,O321,O322,O323,O324,O325,O326,O327,O328,O329,O330,O331,O332,O333,O334,O335,
O336,O337,O338,O339,O340,O341,O342,O343,O344,O345,O346,O347,O348,O349,O350,O351,O352,O353,O354,O355,O356,
O357,O358,O359,O360,O361,O362,O363,O364,O365,O366,O367,O368,O369,O370,O371,O372,O373,O374,O375,O376,O377,
O378,O379,O380,O381,O382,O383,O384,O385,O386,O387,O388,O389,O390,O391,O392,O393,O394,O395,O396,O397,O398,
O399,O400,O401,O402,O403,O404,O405,O406,O407,O408,O409,O410,O411,O412,O413,O414,O415,O416,O417,O418,O419,
O420,O421,O422,O423,O424,O425,O426,O427,O428,O429,O430,O431,O432,O433,O434,O435,O436,O437,O438,O439,O440,
O441,O442,O443,O444,O445,O446,O447,O448,O449,O450,O451,O452,O453,O454,O455,O456,O457,O458,O459,O460,O461,
O462,O463,O464,O465,O466,O467,O468,O469,O470,O471,O472,O473,O474,O475,O476,O477,O478,O479,O480,O481,O482,
O483,O484,O485,O486,O487,O488,O489,O490,O491,O492,O493,O494,O495,O496,O497,O498,O499,O500,O501,O502,O503,
O504,O505,O506,O507,O508,O509,O510,O511,O512,O513,O514,O515,O516,O517,O518,O519,O520,O521,O522,O523,O524,
O525,O526,O527,O528,O529,O530,O531,O532,O533,O534,O535,O536,O537,O538,O539,O540,O541,O542,O543,O544,O545,
O546,O547,O548,O549,O550,O551,O552,O553,O554,O555,O556,O557,O558,O559,O560,O561,O562,O563,O564,O565,O566,
O567,O568,O569,O570,O571,O572,O573,O574,O575,O576,O577,O578,O579,O580,O581,O582,O583,O584,O585,O586,O587,
O588,O589,O590,O591,O592,O593,O594,O595,O596,O597,O598,O599,O600,O601,O602,O603,O604,O605,O606,O607,O608,
O609,O610,O611,O612,O613,O614,O615,O616,O617,O618,O619,O620,O621,O622,O623,O624,O625,O626,O627,O628,O629,
O630,O631,O632,O633,O634,O635,O636,O637,O638,O639,O640,O641,O642,O643,O644,O645,O646,O647,O648,O649,O650,
O651,O652,O653,O654,O655,O656,O657,O658,O659,O660,O661,O662,O663,O664,O665,O666,O667,O668,O669,O670,O671,
O672,O673,O674,O675,O676,O677,O678,O679,O680,O681,O682,O683,O684,O685,O686,O687,O688,O689,O690,O691,O692,
O693,O694,O695,O696,O697,O698,O699,O700,O701,O702,O703,O704,O705,O706,O707,O708,O709,O710,O711,O712,O713,
O714,O715,O716,O717,O718,O719,O720,O721,O722,O723,O724,O725,O726,O727,O728,O729,O730,O731,O732,O733,O734,
O735,O736,O737,O738,O739,O740,O741,O742,O743,O744,O745,O746,O747,O748,O749,O750,O751,O752,O753,O754,O755,
O756,O757,O758,O759,O760,O761,O762,O763,O764,O765,O766,O767,O768,O769,O770,O771,O772,O773,O774,O775,O776,
O777,O778,O779,O780,O781,O782,O783,O784,O785,O786,O787,O788,O789,O790,O791,O792,O793,O794,O795,O796,O797,
O798,O799,O800,O801,O802,O803,O804,O805,O806,O807,O808,O809,O810,O811,O812,O813,O814,O815,O816,O817,O818,
O819,O820,O821,O822,O823,O824,O825,O826,O827,O828,O829,O830,O831,O832,O833,O834,O835,O836,O837,O838,O839,
O840,O841,O842,O843,O844,O845,O846,O847,O848,O849,O850,O851,O852,O853,O854,O855,O856,O857,O858,O859,O860,
O861,O862,O863,O864,O865,O866,O867,O868,O869,O870,O871,O872,O873,O874,O875,O876,O877,O878,O879,O880,O881,
O882,O883,O884,O885,O886,O887,O888,O889,O890,O891,O892,O893,O894,O895,O896,O897,O898,O899,O900,O901,O902,
O903,O904,O905,O906,O907,O908,O909,O910,O911,O912,O913,O914,O915,O916,O917,O918,O919,O920,O921,O922,O923,
O924,O925,O926,O927,O928,O929,O930,O931,O932,O933,O934,O935,O936,O937,O938,O939,O940,O941,O942,O943,O944,
O945,O946,O947,O948,O949,O950,O951,O952,O953,O954,O955,O956,O957,O958,O959,O960,O961,O962,O963,O964,O965,
O966,O967,O968,O969,O970,O971,O972,O973,O974,O975,O976,O977,O978,O979,O980,O981,O982,O983,O984,O985,O986,
O987,O988,O989,O990,O991,O992,O993,O994,O995,O996,O997,O998,O999,O1000,O1001,O1002,O1003,O1004,O1005,O1006,O1007,
O1008,O1009,O1010,O1011,O1012,O1013,O1014,O1015,O1016,O1017,O1018,O1019,O1020,O1021,O1022,O1023,O1024,O1025,O1026,O1027,O1028,
O1029,O1030,O1031,O1032,O1033,O1034,O1035,O1036,O1037,O1038,O1039,O1040,O1041,O1042,O1043,O1044,O1045,O1046,O1047,O1048,O1049,
O1050,O1051,O1052,O1053,O1054,O1055,O1056,O1057,O1058,O1059,O1060,O1061,O1062,O1063,O1064,O1065,O1066,O1067,O1068,O1069,O1070,
O1071,O1072,O1073,O1074,O1075,O1076,O1077,O1078,O1079,O1080,O1081,O1082,O1083,O1084,O1085,O1086,O1087,O1088,O1089,O1090,O1091,
O1092,O1093,O1094,O1095,O1096,O1097,O1098,O1099,O1100,O1101,O1102,O1103,O1104,O1105,O1106,O1107,O1108,O1109,O1110,O1111,O1112,
O1113,O1114,O1115,O1116,O1117,O1118,O1119,O1120,O1121,O1122,O1123,O1124,O1125,O1126,O1127,O1128,O1129,O1130,O1131,O1132,O1133,
O1134,O1135,O1136,O1137,O1138,O1139,O1140,O1141,O1142,O1143,O1144,O1145,O1146,O1147,O1148,O1149,O1150,O1151,O1152,O1153,O1154,
O1155,O1156,O1157,O1158,O1159,O1160,O1161,O1162,O1163,O1164,O1165,O1166,O1167,O1168,O1169,O1170,O1171,O1172,O1173,O1174,O1175,
O1176,O1177,O1178,O1179,O1180,O1181,O1182,O1183,O1184,O1185,O1186,O1187,O1188,O1189,O1190,O1191,O1192,O1193,O1194,O1195,O1196,
O1197,O1198,O1199,O1200,O1201,O1202,O1203,O1204,O1205,O1206,O1207,O1208,O1209,O1210,O1211,O1212,O1213,O1214,O1215,O1216,O1217,
O1218,O1219,O1220,O1221,O1222,O1223,O1224,O1225,O1226,O1227,O1228,O1229,O1230,O1231,O1232,O1233,O1234,O1235,O1236,O1237,O1238,
O1239,O1240,O1241,O1242,O1243,O1244,O1245,O1246,O1247,O1248,O1249,O1250,O1251,O1252,O1253,O1254,O1255,O1256,O1257,O1258,O1259,
O1260,O1261,O1262,O1263,O1264,O1265,O1266,O1267,O1268,O1269,O1270,O1271,O1272,O1273,O1274,O1275,O1276,O1277,O1278,O1279,O1280,
O1281,O1282,O1283,O1284,O1285,O1286,O1287,O1288,O1289,O1290,O1291,O1292,O1293,O1294,O1295,O1296,O1297,O1298,O1299,O1300,O1301,
O1302,O1303,O1304,O1305,O1306,O1307,O1308,O1309,O1310,O1311,O1312,O1313,O1314,O1315,O1316,O1317,O1318,O1319,O1320,O1321,O1322,
O1323,O1324,O1325,O1326,O1327,O1328,O1329,O1330,O1331,O1332,O1333,O1334,O1335,O1336,O1337,O1338,O1339,O1340,O1341,O1342,O1343,
O1344,O1345,O1346,O1347,O1348,O1349,O1350,O1351,O1352,O1353,O1354,O1355,O1356,O1357,O1358,O1359,O1360,O1361,O1362,O1363,O1364,
O1365,O1366,O1367,O1368,O1369,O1370,O1371,O1372,O1373,O1374,O1375,O1376,O1377,O1378,O1379,O1380,O1381,O1382,O1383,O1384,O1385,
O1386,O1387,O1388,O1389,O1390,O1391,O1392,O1393,O1394,O1395,O1396,O1397);
input I1;
input I2;
input I3;
input I4;
input I5;
input I6;
input I7;
input I8;
input I9;
input I10;
input I11;
input I12;
input I13;
input I14;
input I15;
input I16;
input I17;
input I18;
input I19;
input I20;
input I21;
input I22;
input I23;
input I24;
input I25;
input I26;
input I27;
input I28;
input I29;
input I30;
input I31;
input I32;
input I33;
input I34;
input I35;
input I36;
input I37;
input I38;
input I39;
input I40;
input I41;
input I42;
input I43;
input I44;
input I45;
input I46;
input I47;
input I48;
input I49;
input I50;
input I51;
input I52;
input I53;
input I54;
input I55;
input I56;
input I57;
input I58;
input I59;
input I60;
input I61;
input I62;
input I63;
input I64;
input I65;
input I66;
input I67;
input I68;
input I69;
input I70;
input I71;
input I72;
input I73;
input I74;
input I75;
input I76;
input I77;
input I78;
input I79;
input I80;
input I81;
input I82;
input I83;
input I84;
input I85;
input I86;
input I87;
input I88;
input I89;
input I90;
input I91;
input I92;
input I93;
input I94;
input I95;
input I96;
input I97;
input I98;
input I99;
input I100;
input I101;
input I102;
input I103;
input I104;
input I105;
input I106;
input I107;
input I108;
input I109;
input I110;
input I111;
input I112;
input I113;
input I114;
input I115;
input I116;
input I117;
input I118;
input I119;
input I120;
input I121;
input I122;
input I123;
input I124;
input I125;
input I126;
input I127;
input I128;
input I129;
input I130;
input I131;
input I132;
input I133;
input I134;
input I135;
input I136;
input I137;
input I138;
input I139;
input I140;
input I141;
input I142;
input I143;
input I144;
input I145;
input I146;
input I147;
input I148;
input I149;
input I150;
input I151;
input I152;
input I153;
input I154;
input I155;
input I156;
input I157;
input I158;
input I159;
input I160;
input I161;
input I162;
input I163;
input I164;
input I165;
input I166;
input I167;
input I168;
input I169;
input I170;
input I171;
input I172;
input I173;
input I174;
input I175;
input I176;
input I177;
input I178;
input I179;
input I180;
input I181;
input I182;
input I183;
input I184;
input I185;
input I186;
input I187;
input I188;
input I189;
input I190;
input I191;
input I192;
input I193;
input I194;
input I195;
input I196;
input I197;
input I198;
input I199;
input I200;
input I201;
input I202;
input I203;
input I204;
input I205;
input I206;
input I207;
input I208;
input I209;
input I210;
input I211;
input I212;
input I213;
input I214;
input I215;
input I216;
input I217;
input I218;
input I219;
input I220;
input I221;
input I222;
input I223;
input I224;
input I225;
input I226;
input I227;
input I228;
input I229;
input I230;
input I231;
input I232;
input I233;
input I234;
input I235;
input I236;
input I237;
input I238;
input I239;
input I240;
input I241;
input I242;
input I243;
input I244;
input I245;
input I246;
input I247;
input I248;
input I249;
input I250;
input I251;
input I252;
input I253;
input I254;
input I255;
input I256;
input I257;
input I258;
input I259;
input I260;
input I261;
input I262;
input I263;
input I264;
input I265;
input I266;
input I267;
input I268;
input I269;
input I270;
input I271;
input I272;
input I273;
input I274;
input I275;
input I276;
input I277;
input I278;
input I279;
input I280;
input I281;
input I282;
input I283;
input I284;
input I285;
input I286;
input I287;
input I288;
input I289;
input I290;
input I291;
input I292;
input I293;
input I294;
input I295;
input I296;
input I297;
input I298;
input I299;
input I300;
input I301;
input I302;
input I303;
input I304;
input I305;
input I306;
input I307;
input I308;
input I309;
input I310;
input I311;
input I312;
input I313;
input I314;
input I315;
input I316;
input I317;
input I318;
input I319;
input I320;
input I321;
input I322;
input I323;
input I324;
input I325;
input I326;
input I327;
input I328;
input I329;
input I330;
input I331;
input I332;
input I333;
input I334;
input I335;
input I336;
input I337;
input I338;
input I339;
input I340;
input I341;
input I342;
input I343;
input I344;
input I345;
input I346;
input I347;
input I348;
input I349;
input I350;
input I351;
input I352;
input I353;
input I354;
input I355;
input I356;
input I357;
input I358;
input I359;
input I360;
input I361;
input I362;
input I363;
input I364;
input I365;
input I366;
input I367;
input I368;
input I369;
input I370;
input I371;
input I372;
input I373;
input I374;
input I375;
input I376;
input I377;
input I378;
input I379;
input I380;
input I381;
input I382;
input I383;
input I384;
input I385;
input I386;
input I387;
input I388;
input I389;
input I390;
input I391;
input I392;
input I393;
input I394;
input I395;
input I396;
input I397;
input I398;
input I399;
input I400;
input I401;
input I402;
input I403;
input I404;
input I405;
input I406;
input I407;
input I408;
input I409;
input I410;
input I411;
input I412;
input I413;
input I414;
input I415;
input I416;
input I417;
input I418;
input I419;
input I420;
input I421;
input I422;
input I423;
input I424;
input I425;
input I426;
input I427;
input I428;
input I429;
input I430;
input I431;
input I432;
input I433;
input I434;
input I435;
input I436;
input I437;
input I438;
input I439;
input I440;
input I441;
input I442;
input I443;
input I444;
input I445;
input I446;
input I447;
input I448;
input I449;
input I450;
input I451;
input I452;
input I453;
input I454;
input I455;
input I456;
input I457;
input I458;
input I459;
input I460;
input I461;
input I462;
input I463;
input I464;
input I465;
input I466;
input I467;
input I468;
input I469;
input I470;
input I471;
input I472;
input I473;
input I474;
input I475;
input I476;
input I477;
input I478;
input I479;
input I480;
input I481;
input I482;
input I483;
input I484;
input I485;
input I486;
input I487;
input I488;
input I489;
input I490;
input I491;
input I492;
input I493;
input I494;
input I495;
input I496;
input I497;
input I498;
input I499;
input I500;
input I501;
input I502;
input I503;
input I504;
input I505;
input I506;
input I507;
input I508;
input I509;
input I510;
input I511;
input I512;
input I513;
input I514;
input I515;
input I516;
input I517;
input I518;
input I519;
input I520;
input I521;
input I522;
input I523;
input I524;
input I525;
input I526;
input I527;
input I528;
input I529;
input I530;
input I531;
input I532;
input I533;
input I534;
input I535;
input I536;
input I537;
input I538;
input I539;
input I540;
input I541;
input I542;
input I543;
input I544;
input I545;
input I546;
input I547;
input I548;
input I549;
input I550;
input I551;
input I552;
input I553;
input I554;
input I555;
input I556;
input I557;
input I558;
input I559;
input I560;
input I561;
input I562;
input I563;
input I564;
input I565;
input I566;
input I567;
input I568;
input I569;
input I570;
input I571;
input I572;
input I573;
input I574;
input I575;
input I576;
input I577;
input I578;
input I579;
input I580;
input I581;
input I582;
input I583;
input I584;
input I585;
input I586;
input I587;
input I588;
input I589;
input I590;
input I591;
input I592;
input I593;
input I594;
input I595;
input I596;
input I597;
input I598;
input I599;
input I600;
input I601;
input I602;
input I603;
input I604;
input I605;
input I606;
input I607;
input I608;
input I609;
input I610;
input I611;
input I612;
input I613;
input I614;
input I615;
input I616;
input I617;
input I618;
input I619;
input I620;
input I621;
input I622;
input I623;
input I624;
input I625;
input I626;
input I627;
input I628;
input I629;
input I630;
input I631;
input I632;
input I633;
input I634;
input I635;
input I636;
input I637;
input I638;
input I639;
input I640;
input I641;
input I642;
input I643;
input I644;
input I645;
input I646;
input I647;
input I648;
input I649;
input I650;
input I651;
input I652;
input I653;
input I654;
input I655;
input I656;
input I657;
input I658;
input I659;
input I660;
input I661;
input I662;
input I663;
input I664;
input I665;
input I666;
input I667;
input I668;
input I669;
input I670;
input I671;
input I672;
input I673;
input I674;
input I675;
input I676;
input I677;
input I678;
input I679;
input I680;
input I681;
input I682;
input I683;
input I684;
input I685;
input I686;
input I687;
input I688;
input I689;
input I690;
input I691;
input I692;
input I693;
input I694;
input I695;
input I696;
input I697;
input I698;
input I699;
input I700;
input I701;
input I702;
input I703;
input I704;
input I705;
input I706;
input I707;
input I708;
input I709;
input I710;
input I711;
input I712;
input I713;
input I714;
input I715;
input I716;
input I717;
input I718;
input I719;
input I720;
input I721;
input I722;
input I723;
input I724;
input I725;
input I726;
input I727;
input I728;
input I729;
input I730;
input I731;
input I732;
input I733;
input I734;
input I735;
input I736;
input I737;
input I738;
input I739;
input I740;
input I741;
input I742;
input I743;
input I744;
input I745;
input I746;
input I747;
input I748;
input I749;
input I750;
input I751;
input I752;
input I753;
input I754;
input I755;
input I756;
input I757;
input I758;
input I759;
input I760;
input I761;
input I762;
input I763;
input I764;
input I765;
input I766;
input I767;
input I768;
input I769;
input I770;
input I771;
input I772;
input I773;
input I774;
input I775;
input I776;
input I777;
input I778;
input I779;
input I780;
input I781;
input I782;
input I783;
input I784;
input I785;
input I786;
input I787;
input I788;
input I789;
input I790;
input I791;
input I792;
input I793;
input I794;
input I795;
input I796;
input I797;
input I798;
input I799;
input I800;
input I801;
input I802;
input I803;
input I804;
input I805;
input I806;
input I807;
input I808;
input I809;
input I810;
input I811;
input I812;
input I813;
input I814;
input I815;
input I816;
input I817;
input I818;
input I819;
input I820;
input I821;
input I822;
input I823;
input I824;
input I825;
input I826;
input I827;
input I828;
input I829;
input I830;
input I831;
input I832;
input I833;
input I834;
input I835;
input I836;
input I837;
input I838;
input I839;
input I840;
input I841;
input I842;
input I843;
input I844;
input I845;
input I846;
input I847;
input I848;
input I849;
input I850;
input I851;
input I852;
input I853;
input I854;
input I855;
input I856;
input I857;
input I858;
input I859;
input I860;
input I861;
input I862;
input I863;
input I864;
input I865;
input I866;
input I867;
input I868;
input I869;
input I870;
input I871;
input I872;
input I873;
input I874;
input I875;
input I876;
input I877;
input I878;
input I879;
input I880;
input I881;
input I882;
input I883;
input I884;
input I885;
input I886;
input I887;
input I888;
input I889;
input I890;
input I891;
input I892;
input I893;
input I894;
input I895;
input I896;
input I897;
input I898;
input I899;
input I900;
input I901;
input I902;
input I903;
input I904;
input I905;
input I906;
input I907;
input I908;
input I909;
input I910;
input I911;
input I912;
input I913;
input I914;
input I915;
input I916;
input I917;
input I918;
input I919;
input I920;
input I921;
input I922;
input I923;
input I924;
input I925;
input I926;
input I927;
input I928;
input I929;
input I930;
input I931;
input I932;
input I933;
input I934;
input I935;
input I936;
input I937;
input I938;
input I939;
input I940;
input I941;
input I942;
input I943;
input I944;
input I945;
input I946;
input I947;
input I948;
input I949;
input I950;
input I951;
input I952;
input I953;
input I954;
input I955;
input I956;
input I957;
input I958;
input I959;
input I960;
input I961;
input I962;
input I963;
input I964;
input I965;
input I966;
input I967;
input I968;
input I969;
input I970;
input I971;
input I972;
input I973;
input I974;
input I975;
input I976;
input I977;
input I978;
input I979;
input I980;
input I981;
input I982;
input I983;
input I984;
input I985;
input I986;
input I987;
input I988;
input I989;
input I990;
input I991;
input I992;
input I993;
input I994;
input I995;
input I996;
input I997;
input I998;
input I999;
input I1000;
input I1001;
input I1002;
input I1003;
input I1004;
input I1005;
input I1006;
input I1007;
input I1008;
input I1009;
input I1010;
input I1011;
input I1012;
input I1013;
input I1014;
input I1015;
input I1016;
input I1017;
input I1018;
input I1019;
input I1020;
input I1021;
input I1022;
input I1023;
input I1024;
input I1025;
input I1026;
input I1027;
input I1028;
input I1029;
input I1030;
input I1031;
input I1032;
input I1033;
input I1034;
input I1035;
input I1036;
input I1037;
input I1038;
input I1039;
input I1040;
input I1041;
input I1042;
input I1043;
input I1044;
input I1045;
input I1046;
input I1047;
input I1048;
input I1049;
input I1050;
input I1051;
input I1052;
input I1053;
input I1054;
input I1055;
input I1056;
input I1057;
input I1058;
input I1059;
input I1060;
input I1061;
input I1062;
input I1063;
input I1064;
input I1065;
input I1066;
input I1067;
input I1068;
input I1069;
input I1070;
input I1071;
input I1072;
input I1073;
input I1074;
input I1075;
input I1076;
input I1077;
input I1078;
input I1079;
input I1080;
input I1081;
input I1082;
input I1083;
input I1084;
input I1085;
input I1086;
input I1087;
input I1088;
input I1089;
input I1090;
input I1091;
input I1092;
input I1093;
input I1094;
input I1095;
input I1096;
input I1097;
input I1098;
input I1099;
input I1100;
input I1101;
input I1102;
input I1103;
input I1104;
input I1105;
input I1106;
input I1107;
input I1108;
input I1109;
input I1110;
input I1111;
input I1112;
input I1113;
input I1114;
input I1115;
input I1116;
input I1117;
input I1118;
input I1119;
input I1120;
input I1121;
input I1122;
input I1123;
input I1124;
input I1125;
input I1126;
input I1127;
input I1128;
input I1129;
input I1130;
input I1131;
input I1132;
input I1133;
input I1134;
input I1135;
input I1136;
input I1137;
input I1138;
input I1139;
input I1140;
input I1141;
input I1142;
input I1143;
input I1144;
input I1145;
input I1146;
input I1147;
input I1148;
input I1149;
input I1150;
input I1151;
input I1152;
input I1153;
input I1154;
input I1155;
input I1156;
input I1157;
input I1158;
input I1159;
input I1160;
input I1161;
input I1162;
input I1163;
input I1164;
input I1165;
input I1166;
input I1167;
input I1168;
input I1169;
input I1170;
input I1171;
input I1172;
input I1173;
input I1174;
input I1175;
input I1176;
input I1177;
input I1178;
input I1179;
input I1180;
input I1181;
input I1182;
input I1183;
input I1184;
input I1185;
input I1186;
input I1187;
input I1188;
input I1189;
input I1190;
input I1191;
input I1192;
input I1193;
input I1194;
input I1195;
input I1196;
input I1197;
input I1198;
input I1199;
input I1200;
input I1201;
input I1202;
input I1203;
input I1204;
input I1205;
input I1206;
input I1207;
input I1208;
input I1209;
input I1210;
input I1211;
input I1212;
input I1213;
input I1214;
input I1215;
input I1216;
input I1217;
input I1218;
input I1219;
input I1220;
input I1221;
input I1222;
input I1223;
input I1224;
input I1225;
input I1226;
input I1227;
input I1228;
input I1229;
input I1230;
input I1231;
input I1232;
input I1233;
input I1234;
input I1235;
input I1236;
input I1237;
input I1238;
input I1239;
input I1240;
input I1241;
input I1242;
input I1243;
input I1244;
input I1245;
input I1246;
input I1247;
input I1248;
input I1249;
input I1250;
input I1251;
input I1252;
input I1253;
input I1254;
input I1255;
input I1256;
input I1257;
input I1258;
input I1259;
input I1260;
input I1261;
input I1262;
input I1263;
input I1264;
input I1265;
input I1266;
input I1267;
input I1268;
input I1269;
input I1270;
input I1271;
input I1272;
input I1273;
input I1274;
input I1275;
input I1276;
input I1277;
input I1278;
input I1279;
input I1280;
input I1281;
input I1282;
input I1283;
input I1284;
input I1285;
input I1286;
input I1287;
input I1288;
input I1289;
input I1290;
input I1291;
input I1292;
input I1293;
input I1294;
input I1295;
input I1296;
input I1297;
input I1298;
input I1299;
input I1300;
input I1301;
input I1302;
input I1303;
input I1304;
input I1305;
input I1306;
input I1307;
input I1308;
input I1309;
input I1310;
input I1311;
input I1312;
input I1313;
input I1314;
input I1315;
input I1316;
input I1317;
input I1318;
input I1319;
input I1320;
input I1321;
input I1322;
input I1323;
input I1324;
input I1325;
input I1326;
input I1327;
input I1328;
input I1329;
input I1330;
input I1331;
input I1332;
input I1333;
input I1334;
input I1335;
input I1336;
input I1337;
input I1338;
input I1339;
input I1340;
input I1341;
input I1342;
input I1343;
input I1344;
input I1345;
input I1346;
input I1347;
input I1348;
input I1349;
input I1350;
input I1351;
input I1352;
input I1353;
input I1354;
input I1355;
input I1356;
input I1357;
input I1358;
input I1359;
input I1360;
input I1361;
input I1362;
input I1363;
input I1364;
input I1365;
input I1366;
input I1367;
input I1368;
input I1369;
input I1370;
input I1371;
input I1372;
input I1373;
input I1374;
input I1375;
input I1376;
input I1377;
input I1378;
input I1379;
input I1380;
input I1381;
input I1382;
input I1383;
input I1384;
input I1385;
input I1386;
input I1387;
input I1388;
input I1389;
input I1390;
input I1391;
input I1392;
input I1393;
input I1394;
input I1395;
input I1396;
input I1397;
input I1398;
input I1399;
input I1400;
input I1401;
input I1402;
input I1403;
input I1404;
input I1405;
input I1406;
input I1407;
input I1408;
input I1409;
input I1410;
input I1411;
input I1412;
input I1413;
input I1414;
input I1415;
input I1416;
input I1417;
input I1418;
input I1419;
input I1420;
input I1421;
input I1422;
input I1423;
input I1424;
input I1425;
input I1426;
input I1427;
input I1428;
input I1429;
input I1430;
input I1431;
input I1432;
input I1433;
input I1434;
input I1435;
input I1436;
input I1437;
input I1438;
input I1439;
input I1440;
input I1441;
input I1442;
input I1443;
input I1444;
input I1445;
input I1446;
input I1447;
input I1448;
input I1449;
input I1450;
input I1451;
input I1452;
input I1453;
input I1454;
input I1455;
input I1456;
input I1457;
input I1458;
input I1459;
input I1460;
input I1461;
input I1462;
input I1463;
input I1464;
input I1465;
input I1466;
input I1467;
input I1468;
input I1469;
input I1470;
input I1471;
input I1472;
input I1473;
input I1474;
input I1475;
input I1476;
input I1477;
input I1478;
input I1479;
input I1480;
input I1481;
input I1482;
input I1483;
input I1484;
input I1485;
input I1486;
input I1487;
input I1488;
input I1489;
input I1490;
input I1491;
input I1492;
input I1493;
input I1494;
input I1495;
input I1496;
input I1497;
input I1498;
input I1499;
input I1500;
input I1501;
input I1502;
input I1503;
input I1504;
input I1505;
input I1506;
input I1507;
input I1508;
input I1509;
input I1510;
input I1511;
input I1512;
input I1513;
input I1514;
input I1515;
input I1516;
input I1517;
input I1518;
input I1519;
input I1520;
input I1521;
input I1522;
input I1523;
input I1524;
input I1525;
input I1526;
input I1527;
input I1528;
input I1529;
input I1530;
input I1531;
input I1532;
input I1533;
input I1534;
input I1535;
input I1536;
input I1537;
input I1538;
input I1539;
input I1540;
input I1541;
input I1542;
input I1543;
input I1544;
input I1545;
input I1546;
input I1547;
input I1548;
input I1549;
input I1550;
input I1551;
input I1552;
input I1553;
input I1554;
input I1555;
input I1556;
input I1557;
input I1558;
input I1559;
input I1560;
input I1561;
input I1562;
input I1563;
input I1564;
input I1565;
input I1566;
input I1567;
input I1568;
input I1569;
input I1570;
input I1571;
input I1572;
input I1573;
input I1574;
input I1575;
input I1576;
input I1577;
input I1578;
input I1579;
input I1580;
input I1581;
input I1582;
input I1583;
input I1584;
input I1585;
input I1586;
input I1587;
input I1588;
input I1589;
input I1590;
input I1591;
input I1592;
input I1593;
input I1594;
input I1595;
input I1596;
input I1597;
input I1598;
input I1599;
input I1600;
input I1601;
input I1602;
input I1603;
input I1604;
input I1605;
input I1606;
input I1607;
input I1608;
input I1609;
input I1610;
input I1611;
input I1612;
input I1613;
input I1614;
input I1615;
input I1616;
input I1617;
input I1618;
input I1619;
input I1620;
input I1621;
input I1622;
input I1623;
input I1624;
input I1625;
input I1626;
input I1627;
input I1628;
input I1629;
input I1630;
input I1631;
input I1632;
input I1633;
input I1634;
input I1635;
input I1636;
input I1637;
input I1638;
input I1639;
input I1640;
input I1641;
input I1642;
input I1643;
input I1644;

output O1;
output O2;
output O3;
output O4;
output O5;
output O6;
output O7;
output O8;
output O9;
output O10;
output O11;
output O12;
output O13;
output O14;
output O15;
output O16;
output O17;
output O18;
output O19;
output O20;
output O21;
output O22;
output O23;
output O24;
output O25;
output O26;
output O27;
output O28;
output O29;
output O30;
output O31;
output O32;
output O33;
output O34;
output O35;
output O36;
output O37;
output O38;
output O39;
output O40;
output O41;
output O42;
output O43;
output O44;
output O45;
output O46;
output O47;
output O48;
output O49;
output O50;
output O51;
output O52;
output O53;
output O54;
output O55;
output O56;
output O57;
output O58;
output O59;
output O60;
output O61;
output O62;
output O63;
output O64;
output O65;
output O66;
output O67;
output O68;
output O69;
output O70;
output O71;
output O72;
output O73;
output O74;
output O75;
output O76;
output O77;
output O78;
output O79;
output O80;
output O81;
output O82;
output O83;
output O84;
output O85;
output O86;
output O87;
output O88;
output O89;
output O90;
output O91;
output O92;
output O93;
output O94;
output O95;
output O96;
output O97;
output O98;
output O99;
output O100;
output O101;
output O102;
output O103;
output O104;
output O105;
output O106;
output O107;
output O108;
output O109;
output O110;
output O111;
output O112;
output O113;
output O114;
output O115;
output O116;
output O117;
output O118;
output O119;
output O120;
output O121;
output O122;
output O123;
output O124;
output O125;
output O126;
output O127;
output O128;
output O129;
output O130;
output O131;
output O132;
output O133;
output O134;
output O135;
output O136;
output O137;
output O138;
output O139;
output O140;
output O141;
output O142;
output O143;
output O144;
output O145;
output O146;
output O147;
output O148;
output O149;
output O150;
output O151;
output O152;
output O153;
output O154;
output O155;
output O156;
output O157;
output O158;
output O159;
output O160;
output O161;
output O162;
output O163;
output O164;
output O165;
output O166;
output O167;
output O168;
output O169;
output O170;
output O171;
output O172;
output O173;
output O174;
output O175;
output O176;
output O177;
output O178;
output O179;
output O180;
output O181;
output O182;
output O183;
output O184;
output O185;
output O186;
output O187;
output O188;
output O189;
output O190;
output O191;
output O192;
output O193;
output O194;
output O195;
output O196;
output O197;
output O198;
output O199;
output O200;
output O201;
output O202;
output O203;
output O204;
output O205;
output O206;
output O207;
output O208;
output O209;
output O210;
output O211;
output O212;
output O213;
output O214;
output O215;
output O216;
output O217;
output O218;
output O219;
output O220;
output O221;
output O222;
output O223;
output O224;
output O225;
output O226;
output O227;
output O228;
output O229;
output O230;
output O231;
output O232;
output O233;
output O234;
output O235;
output O236;
output O237;
output O238;
output O239;
output O240;
output O241;
output O242;
output O243;
output O244;
output O245;
output O246;
output O247;
output O248;
output O249;
output O250;
output O251;
output O252;
output O253;
output O254;
output O255;
output O256;
output O257;
output O258;
output O259;
output O260;
output O261;
output O262;
output O263;
output O264;
output O265;
output O266;
output O267;
output O268;
output O269;
output O270;
output O271;
output O272;
output O273;
output O274;
output O275;
output O276;
output O277;
output O278;
output O279;
output O280;
output O281;
output O282;
output O283;
output O284;
output O285;
output O286;
output O287;
output O288;
output O289;
output O290;
output O291;
output O292;
output O293;
output O294;
output O295;
output O296;
output O297;
output O298;
output O299;
output O300;
output O301;
output O302;
output O303;
output O304;
output O305;
output O306;
output O307;
output O308;
output O309;
output O310;
output O311;
output O312;
output O313;
output O314;
output O315;
output O316;
output O317;
output O318;
output O319;
output O320;
output O321;
output O322;
output O323;
output O324;
output O325;
output O326;
output O327;
output O328;
output O329;
output O330;
output O331;
output O332;
output O333;
output O334;
output O335;
output O336;
output O337;
output O338;
output O339;
output O340;
output O341;
output O342;
output O343;
output O344;
output O345;
output O346;
output O347;
output O348;
output O349;
output O350;
output O351;
output O352;
output O353;
output O354;
output O355;
output O356;
output O357;
output O358;
output O359;
output O360;
output O361;
output O362;
output O363;
output O364;
output O365;
output O366;
output O367;
output O368;
output O369;
output O370;
output O371;
output O372;
output O373;
output O374;
output O375;
output O376;
output O377;
output O378;
output O379;
output O380;
output O381;
output O382;
output O383;
output O384;
output O385;
output O386;
output O387;
output O388;
output O389;
output O390;
output O391;
output O392;
output O393;
output O394;
output O395;
output O396;
output O397;
output O398;
output O399;
output O400;
output O401;
output O402;
output O403;
output O404;
output O405;
output O406;
output O407;
output O408;
output O409;
output O410;
output O411;
output O412;
output O413;
output O414;
output O415;
output O416;
output O417;
output O418;
output O419;
output O420;
output O421;
output O422;
output O423;
output O424;
output O425;
output O426;
output O427;
output O428;
output O429;
output O430;
output O431;
output O432;
output O433;
output O434;
output O435;
output O436;
output O437;
output O438;
output O439;
output O440;
output O441;
output O442;
output O443;
output O444;
output O445;
output O446;
output O447;
output O448;
output O449;
output O450;
output O451;
output O452;
output O453;
output O454;
output O455;
output O456;
output O457;
output O458;
output O459;
output O460;
output O461;
output O462;
output O463;
output O464;
output O465;
output O466;
output O467;
output O468;
output O469;
output O470;
output O471;
output O472;
output O473;
output O474;
output O475;
output O476;
output O477;
output O478;
output O479;
output O480;
output O481;
output O482;
output O483;
output O484;
output O485;
output O486;
output O487;
output O488;
output O489;
output O490;
output O491;
output O492;
output O493;
output O494;
output O495;
output O496;
output O497;
output O498;
output O499;
output O500;
output O501;
output O502;
output O503;
output O504;
output O505;
output O506;
output O507;
output O508;
output O509;
output O510;
output O511;
output O512;
output O513;
output O514;
output O515;
output O516;
output O517;
output O518;
output O519;
output O520;
output O521;
output O522;
output O523;
output O524;
output O525;
output O526;
output O527;
output O528;
output O529;
output O530;
output O531;
output O532;
output O533;
output O534;
output O535;
output O536;
output O537;
output O538;
output O539;
output O540;
output O541;
output O542;
output O543;
output O544;
output O545;
output O546;
output O547;
output O548;
output O549;
output O550;
output O551;
output O552;
output O553;
output O554;
output O555;
output O556;
output O557;
output O558;
output O559;
output O560;
output O561;
output O562;
output O563;
output O564;
output O565;
output O566;
output O567;
output O568;
output O569;
output O570;
output O571;
output O572;
output O573;
output O574;
output O575;
output O576;
output O577;
output O578;
output O579;
output O580;
output O581;
output O582;
output O583;
output O584;
output O585;
output O586;
output O587;
output O588;
output O589;
output O590;
output O591;
output O592;
output O593;
output O594;
output O595;
output O596;
output O597;
output O598;
output O599;
output O600;
output O601;
output O602;
output O603;
output O604;
output O605;
output O606;
output O607;
output O608;
output O609;
output O610;
output O611;
output O612;
output O613;
output O614;
output O615;
output O616;
output O617;
output O618;
output O619;
output O620;
output O621;
output O622;
output O623;
output O624;
output O625;
output O626;
output O627;
output O628;
output O629;
output O630;
output O631;
output O632;
output O633;
output O634;
output O635;
output O636;
output O637;
output O638;
output O639;
output O640;
output O641;
output O642;
output O643;
output O644;
output O645;
output O646;
output O647;
output O648;
output O649;
output O650;
output O651;
output O652;
output O653;
output O654;
output O655;
output O656;
output O657;
output O658;
output O659;
output O660;
output O661;
output O662;
output O663;
output O664;
output O665;
output O666;
output O667;
output O668;
output O669;
output O670;
output O671;
output O672;
output O673;
output O674;
output O675;
output O676;
output O677;
output O678;
output O679;
output O680;
output O681;
output O682;
output O683;
output O684;
output O685;
output O686;
output O687;
output O688;
output O689;
output O690;
output O691;
output O692;
output O693;
output O694;
output O695;
output O696;
output O697;
output O698;
output O699;
output O700;
output O701;
output O702;
output O703;
output O704;
output O705;
output O706;
output O707;
output O708;
output O709;
output O710;
output O711;
output O712;
output O713;
output O714;
output O715;
output O716;
output O717;
output O718;
output O719;
output O720;
output O721;
output O722;
output O723;
output O724;
output O725;
output O726;
output O727;
output O728;
output O729;
output O730;
output O731;
output O732;
output O733;
output O734;
output O735;
output O736;
output O737;
output O738;
output O739;
output O740;
output O741;
output O742;
output O743;
output O744;
output O745;
output O746;
output O747;
output O748;
output O749;
output O750;
output O751;
output O752;
output O753;
output O754;
output O755;
output O756;
output O757;
output O758;
output O759;
output O760;
output O761;
output O762;
output O763;
output O764;
output O765;
output O766;
output O767;
output O768;
output O769;
output O770;
output O771;
output O772;
output O773;
output O774;
output O775;
output O776;
output O777;
output O778;
output O779;
output O780;
output O781;
output O782;
output O783;
output O784;
output O785;
output O786;
output O787;
output O788;
output O789;
output O790;
output O791;
output O792;
output O793;
output O794;
output O795;
output O796;
output O797;
output O798;
output O799;
output O800;
output O801;
output O802;
output O803;
output O804;
output O805;
output O806;
output O807;
output O808;
output O809;
output O810;
output O811;
output O812;
output O813;
output O814;
output O815;
output O816;
output O817;
output O818;
output O819;
output O820;
output O821;
output O822;
output O823;
output O824;
output O825;
output O826;
output O827;
output O828;
output O829;
output O830;
output O831;
output O832;
output O833;
output O834;
output O835;
output O836;
output O837;
output O838;
output O839;
output O840;
output O841;
output O842;
output O843;
output O844;
output O845;
output O846;
output O847;
output O848;
output O849;
output O850;
output O851;
output O852;
output O853;
output O854;
output O855;
output O856;
output O857;
output O858;
output O859;
output O860;
output O861;
output O862;
output O863;
output O864;
output O865;
output O866;
output O867;
output O868;
output O869;
output O870;
output O871;
output O872;
output O873;
output O874;
output O875;
output O876;
output O877;
output O878;
output O879;
output O880;
output O881;
output O882;
output O883;
output O884;
output O885;
output O886;
output O887;
output O888;
output O889;
output O890;
output O891;
output O892;
output O893;
output O894;
output O895;
output O896;
output O897;
output O898;
output O899;
output O900;
output O901;
output O902;
output O903;
output O904;
output O905;
output O906;
output O907;
output O908;
output O909;
output O910;
output O911;
output O912;
output O913;
output O914;
output O915;
output O916;
output O917;
output O918;
output O919;
output O920;
output O921;
output O922;
output O923;
output O924;
output O925;
output O926;
output O927;
output O928;
output O929;
output O930;
output O931;
output O932;
output O933;
output O934;
output O935;
output O936;
output O937;
output O938;
output O939;
output O940;
output O941;
output O942;
output O943;
output O944;
output O945;
output O946;
output O947;
output O948;
output O949;
output O950;
output O951;
output O952;
output O953;
output O954;
output O955;
output O956;
output O957;
output O958;
output O959;
output O960;
output O961;
output O962;
output O963;
output O964;
output O965;
output O966;
output O967;
output O968;
output O969;
output O970;
output O971;
output O972;
output O973;
output O974;
output O975;
output O976;
output O977;
output O978;
output O979;
output O980;
output O981;
output O982;
output O983;
output O984;
output O985;
output O986;
output O987;
output O988;
output O989;
output O990;
output O991;
output O992;
output O993;
output O994;
output O995;
output O996;
output O997;
output O998;
output O999;
output O1000;
output O1001;
output O1002;
output O1003;
output O1004;
output O1005;
output O1006;
output O1007;
output O1008;
output O1009;
output O1010;
output O1011;
output O1012;
output O1013;
output O1014;
output O1015;
output O1016;
output O1017;
output O1018;
output O1019;
output O1020;
output O1021;
output O1022;
output O1023;
output O1024;
output O1025;
output O1026;
output O1027;
output O1028;
output O1029;
output O1030;
output O1031;
output O1032;
output O1033;
output O1034;
output O1035;
output O1036;
output O1037;
output O1038;
output O1039;
output O1040;
output O1041;
output O1042;
output O1043;
output O1044;
output O1045;
output O1046;
output O1047;
output O1048;
output O1049;
output O1050;
output O1051;
output O1052;
output O1053;
output O1054;
output O1055;
output O1056;
output O1057;
output O1058;
output O1059;
output O1060;
output O1061;
output O1062;
output O1063;
output O1064;
output O1065;
output O1066;
output O1067;
output O1068;
output O1069;
output O1070;
output O1071;
output O1072;
output O1073;
output O1074;
output O1075;
output O1076;
output O1077;
output O1078;
output O1079;
output O1080;
output O1081;
output O1082;
output O1083;
output O1084;
output O1085;
output O1086;
output O1087;
output O1088;
output O1089;
output O1090;
output O1091;
output O1092;
output O1093;
output O1094;
output O1095;
output O1096;
output O1097;
output O1098;
output O1099;
output O1100;
output O1101;
output O1102;
output O1103;
output O1104;
output O1105;
output O1106;
output O1107;
output O1108;
output O1109;
output O1110;
output O1111;
output O1112;
output O1113;
output O1114;
output O1115;
output O1116;
output O1117;
output O1118;
output O1119;
output O1120;
output O1121;
output O1122;
output O1123;
output O1124;
output O1125;
output O1126;
output O1127;
output O1128;
output O1129;
output O1130;
output O1131;
output O1132;
output O1133;
output O1134;
output O1135;
output O1136;
output O1137;
output O1138;
output O1139;
output O1140;
output O1141;
output O1142;
output O1143;
output O1144;
output O1145;
output O1146;
output O1147;
output O1148;
output O1149;
output O1150;
output O1151;
output O1152;
output O1153;
output O1154;
output O1155;
output O1156;
output O1157;
output O1158;
output O1159;
output O1160;
output O1161;
output O1162;
output O1163;
output O1164;
output O1165;
output O1166;
output O1167;
output O1168;
output O1169;
output O1170;
output O1171;
output O1172;
output O1173;
output O1174;
output O1175;
output O1176;
output O1177;
output O1178;
output O1179;
output O1180;
output O1181;
output O1182;
output O1183;
output O1184;
output O1185;
output O1186;
output O1187;
output O1188;
output O1189;
output O1190;
output O1191;
output O1192;
output O1193;
output O1194;
output O1195;
output O1196;
output O1197;
output O1198;
output O1199;
output O1200;
output O1201;
output O1202;
output O1203;
output O1204;
output O1205;
output O1206;
output O1207;
output O1208;
output O1209;
output O1210;
output O1211;
output O1212;
output O1213;
output O1214;
output O1215;
output O1216;
output O1217;
output O1218;
output O1219;
output O1220;
output O1221;
output O1222;
output O1223;
output O1224;
output O1225;
output O1226;
output O1227;
output O1228;
output O1229;
output O1230;
output O1231;
output O1232;
output O1233;
output O1234;
output O1235;
output O1236;
output O1237;
output O1238;
output O1239;
output O1240;
output O1241;
output O1242;
output O1243;
output O1244;
output O1245;
output O1246;
output O1247;
output O1248;
output O1249;
output O1250;
output O1251;
output O1252;
output O1253;
output O1254;
output O1255;
output O1256;
output O1257;
output O1258;
output O1259;
output O1260;
output O1261;
output O1262;
output O1263;
output O1264;
output O1265;
output O1266;
output O1267;
output O1268;
output O1269;
output O1270;
output O1271;
output O1272;
output O1273;
output O1274;
output O1275;
output O1276;
output O1277;
output O1278;
output O1279;
output O1280;
output O1281;
output O1282;
output O1283;
output O1284;
output O1285;
output O1286;
output O1287;
output O1288;
output O1289;
output O1290;
output O1291;
output O1292;
output O1293;
output O1294;
output O1295;
output O1296;
output O1297;
output O1298;
output O1299;
output O1300;
output O1301;
output O1302;
output O1303;
output O1304;
output O1305;
output O1306;
output O1307;
output O1308;
output O1309;
output O1310;
output O1311;
output O1312;
output O1313;
output O1314;
output O1315;
output O1316;
output O1317;
output O1318;
output O1319;
output O1320;
output O1321;
output O1322;
output O1323;
output O1324;
output O1325;
output O1326;
output O1327;
output O1328;
output O1329;
output O1330;
output O1331;
output O1332;
output O1333;
output O1334;
output O1335;
output O1336;
output O1337;
output O1338;
output O1339;
output O1340;
output O1341;
output O1342;
output O1343;
output O1344;
output O1345;
output O1346;
output O1347;
output O1348;
output O1349;
output O1350;
output O1351;
output O1352;
output O1353;
output O1354;
output O1355;
output O1356;
output O1357;
output O1358;
output O1359;
output O1360;
output O1361;
output O1362;
output O1363;
output O1364;
output O1365;
output O1366;
output O1367;
output O1368;
output O1369;
output O1370;
output O1371;
output O1372;
output O1373;
output O1374;
output O1375;
output O1376;
output O1377;
output O1378;
output O1379;
output O1380;
output O1381;
output O1382;
output O1383;
output O1384;
output O1385;
output O1386;
output O1387;
output O1388;
output O1389;
output O1390;
output O1391;
output O1392;
output O1393;
output O1394;
output O1395;
output O1396;
output O1397;

wire W1;
wire W2;
wire W3;
wire W4;
wire W5;
wire W6;
wire W7;
wire W8;
wire W9;
wire W10;
wire W11;
wire W12;
wire W13;
wire W14;
wire W15;
wire W16;
wire W17;
wire W18;
wire W19;
wire W20;
wire W21;
wire W22;
wire W23;
wire W24;
wire W25;
wire W26;
wire W27;
wire W28;
wire W29;
wire W30;
wire W31;
wire W32;
wire W33;
wire W34;
wire W35;
wire W36;
wire W37;
wire W38;
wire W39;
wire W40;
wire W41;
wire W42;
wire W43;
wire W44;
wire W45;
wire W46;
wire W47;
wire W48;
wire W49;
wire W50;
wire W51;
wire W52;
wire W53;
wire W54;
wire W55;
wire W56;
wire W57;
wire W58;
wire W59;
wire W60;
wire W61;
wire W62;
wire W63;
wire W64;
wire W65;
wire W66;
wire W67;
wire W68;
wire W69;
wire W70;
wire W71;
wire W72;
wire W73;
wire W74;
wire W75;
wire W76;
wire W77;
wire W78;
wire W79;
wire W80;
wire W81;
wire W82;
wire W83;
wire W84;
wire W85;
wire W86;
wire W87;
wire W88;
wire W89;
wire W90;
wire W91;
wire W92;
wire W93;
wire W94;
wire W95;
wire W96;
wire W97;
wire W98;
wire W99;
wire W100;
wire W101;
wire W102;
wire W103;
wire W104;
wire W105;
wire W106;
wire W107;
wire W108;
wire W109;
wire W110;
wire W111;
wire W112;
wire W113;
wire W114;
wire W115;
wire W116;
wire W117;
wire W118;
wire W119;
wire W120;
wire W121;
wire W122;
wire W123;
wire W124;
wire W125;
wire W126;
wire W127;
wire W128;
wire W129;
wire W130;
wire W131;
wire W132;
wire W133;
wire W134;
wire W135;
wire W136;
wire W137;
wire W138;
wire W139;
wire W140;
wire W141;
wire W142;
wire W143;
wire W144;
wire W145;
wire W146;
wire W147;
wire W148;
wire W149;
wire W150;
wire W151;
wire W152;
wire W153;
wire W154;
wire W155;
wire W156;
wire W157;
wire W158;
wire W159;
wire W160;
wire W161;
wire W162;
wire W163;
wire W164;
wire W165;
wire W166;
wire W167;
wire W168;
wire W169;
wire W170;
wire W171;
wire W172;
wire W173;
wire W174;
wire W175;
wire W176;
wire W177;
wire W178;
wire W179;
wire W180;
wire W181;
wire W182;
wire W183;
wire W184;
wire W185;
wire W186;
wire W187;
wire W188;
wire W189;
wire W190;
wire W191;
wire W192;
wire W193;
wire W194;
wire W195;
wire W196;
wire W197;
wire W198;
wire W199;
wire W200;
wire W201;
wire W202;
wire W203;
wire W204;
wire W205;
wire W206;
wire W207;
wire W208;
wire W209;
wire W210;
wire W211;
wire W212;
wire W213;
wire W214;
wire W215;
wire W216;
wire W217;
wire W218;
wire W219;
wire W220;
wire W221;
wire W222;
wire W223;
wire W224;
wire W225;
wire W226;
wire W227;
wire W228;
wire W229;
wire W230;
wire W231;
wire W232;
wire W233;
wire W234;
wire W235;
wire W236;
wire W237;
wire W238;
wire W239;
wire W240;
wire W241;
wire W242;
wire W243;
wire W244;
wire W245;
wire W246;
wire W247;
wire W248;
wire W249;
wire W250;
wire W251;
wire W252;
wire W253;
wire W254;
wire W255;
wire W256;
wire W257;
wire W258;
wire W259;
wire W260;
wire W261;
wire W262;
wire W263;
wire W264;
wire W265;
wire W266;
wire W267;
wire W268;
wire W269;
wire W270;
wire W271;
wire W272;
wire W273;
wire W274;
wire W275;
wire W276;
wire W277;
wire W278;
wire W279;
wire W280;
wire W281;
wire W282;
wire W283;
wire W284;
wire W285;
wire W286;
wire W287;
wire W288;
wire W289;
wire W290;
wire W291;
wire W292;
wire W293;
wire W294;
wire W295;
wire W296;
wire W297;
wire W298;
wire W299;
wire W300;
wire W301;
wire W302;
wire W303;
wire W304;
wire W305;
wire W306;
wire W307;
wire W308;
wire W309;
wire W310;
wire W311;
wire W312;
wire W313;
wire W314;
wire W315;
wire W316;
wire W317;
wire W318;
wire W319;
wire W320;
wire W321;
wire W322;
wire W323;
wire W324;
wire W325;
wire W326;
wire W327;
wire W328;
wire W329;
wire W330;
wire W331;
wire W332;
wire W333;
wire W334;
wire W335;
wire W336;
wire W337;
wire W338;
wire W339;
wire W340;
wire W341;
wire W342;
wire W343;
wire W344;
wire W345;
wire W346;
wire W347;
wire W348;
wire W349;
wire W350;
wire W351;
wire W352;
wire W353;
wire W354;
wire W355;
wire W356;
wire W357;
wire W358;
wire W359;
wire W360;
wire W361;
wire W362;
wire W363;
wire W364;
wire W365;
wire W366;
wire W367;
wire W368;
wire W369;
wire W370;
wire W371;
wire W372;
wire W373;
wire W374;
wire W375;
wire W376;
wire W377;
wire W378;
wire W379;
wire W380;
wire W381;
wire W382;
wire W383;
wire W384;
wire W385;
wire W386;
wire W387;
wire W388;
wire W389;
wire W390;
wire W391;
wire W392;
wire W393;
wire W394;
wire W395;
wire W396;
wire W397;
wire W398;
wire W399;
wire W400;
wire W401;
wire W402;
wire W403;
wire W404;
wire W405;
wire W406;
wire W407;
wire W408;
wire W409;
wire W410;
wire W411;
wire W412;
wire W413;
wire W414;
wire W415;
wire W416;
wire W417;
wire W418;
wire W419;
wire W420;
wire W421;
wire W422;
wire W423;
wire W424;
wire W425;
wire W426;
wire W427;
wire W428;
wire W429;
wire W430;
wire W431;
wire W432;
wire W433;
wire W434;
wire W435;
wire W436;
wire W437;
wire W438;
wire W439;
wire W440;
wire W441;
wire W442;
wire W443;
wire W444;
wire W445;
wire W446;
wire W447;
wire W448;
wire W449;
wire W450;
wire W451;
wire W452;
wire W453;
wire W454;
wire W455;
wire W456;
wire W457;
wire W458;
wire W459;
wire W460;
wire W461;
wire W462;
wire W463;
wire W464;
wire W465;
wire W466;
wire W467;
wire W468;
wire W469;
wire W470;
wire W471;
wire W472;
wire W473;
wire W474;
wire W475;
wire W476;
wire W477;
wire W478;
wire W479;
wire W480;
wire W481;
wire W482;
wire W483;
wire W484;
wire W485;
wire W486;
wire W487;
wire W488;
wire W489;
wire W490;
wire W491;
wire W492;
wire W493;
wire W494;
wire W495;
wire W496;
wire W497;
wire W498;
wire W499;
wire W500;
wire W501;
wire W502;
wire W503;
wire W504;
wire W505;
wire W506;
wire W507;
wire W508;
wire W509;
wire W510;
wire W511;
wire W512;
wire W513;
wire W514;
wire W515;
wire W516;
wire W517;
wire W518;
wire W519;
wire W520;
wire W521;
wire W522;
wire W523;
wire W524;
wire W525;
wire W526;
wire W527;
wire W528;
wire W529;
wire W530;
wire W531;
wire W532;
wire W533;
wire W534;
wire W535;
wire W536;
wire W537;
wire W538;
wire W539;
wire W540;
wire W541;
wire W542;
wire W543;
wire W544;
wire W545;
wire W546;
wire W547;
wire W548;
wire W549;
wire W550;
wire W551;
wire W552;
wire W553;
wire W554;
wire W555;
wire W556;
wire W557;
wire W558;
wire W559;
wire W560;
wire W561;
wire W562;
wire W563;
wire W564;
wire W565;
wire W566;
wire W567;
wire W568;
wire W569;
wire W570;
wire W571;
wire W572;
wire W573;
wire W574;
wire W575;
wire W576;
wire W577;
wire W578;
wire W579;
wire W580;
wire W581;
wire W582;
wire W583;
wire W584;
wire W585;
wire W586;
wire W587;
wire W588;
wire W589;
wire W590;
wire W591;
wire W592;
wire W593;
wire W594;
wire W595;
wire W596;
wire W597;
wire W598;
wire W599;
wire W600;
wire W601;
wire W602;
wire W603;
wire W604;
wire W605;
wire W606;
wire W607;
wire W608;
wire W609;
wire W610;
wire W611;
wire W612;
wire W613;
wire W614;
wire W615;
wire W616;
wire W617;
wire W618;
wire W619;
wire W620;
wire W621;
wire W622;
wire W623;
wire W624;
wire W625;
wire W626;
wire W627;
wire W628;
wire W629;
wire W630;
wire W631;
wire W632;
wire W633;
wire W634;
wire W635;
wire W636;
wire W637;
wire W638;
wire W639;
wire W640;
wire W641;
wire W642;
wire W643;
wire W644;
wire W645;
wire W646;
wire W647;
wire W648;
wire W649;
wire W650;
wire W651;
wire W652;
wire W653;
wire W654;
wire W655;
wire W656;
wire W657;
wire W658;
wire W659;
wire W660;
wire W661;
wire W662;
wire W663;
wire W664;
wire W665;
wire W666;
wire W667;
wire W668;
wire W669;
wire W670;
wire W671;
wire W672;
wire W673;
wire W674;
wire W675;
wire W676;
wire W677;
wire W678;
wire W679;
wire W680;
wire W681;
wire W682;
wire W683;
wire W684;
wire W685;
wire W686;
wire W687;
wire W688;
wire W689;
wire W690;
wire W691;
wire W692;
wire W693;
wire W694;
wire W695;
wire W696;
wire W697;
wire W698;
wire W699;
wire W700;
wire W701;
wire W702;
wire W703;
wire W704;
wire W705;
wire W706;
wire W707;
wire W708;
wire W709;
wire W710;
wire W711;
wire W712;
wire W713;
wire W714;
wire W715;
wire W716;
wire W717;
wire W718;
wire W719;
wire W720;
wire W721;
wire W722;
wire W723;
wire W724;
wire W725;
wire W726;
wire W727;
wire W728;
wire W729;
wire W730;
wire W731;
wire W732;
wire W733;
wire W734;
wire W735;
wire W736;
wire W737;
wire W738;
wire W739;
wire W740;
wire W741;
wire W742;
wire W743;
wire W744;
wire W745;
wire W746;
wire W747;
wire W748;
wire W749;
wire W750;
wire W751;
wire W752;
wire W753;
wire W754;
wire W755;
wire W756;
wire W757;
wire W758;
wire W759;
wire W760;
wire W761;
wire W762;
wire W763;
wire W764;
wire W765;
wire W766;
wire W767;
wire W768;
wire W769;
wire W770;
wire W771;
wire W772;
wire W773;
wire W774;
wire W775;
wire W776;
wire W777;
wire W778;
wire W779;
wire W780;
wire W781;
wire W782;
wire W783;
wire W784;
wire W785;
wire W786;
wire W787;
wire W788;
wire W789;
wire W790;
wire W791;
wire W792;
wire W793;
wire W794;
wire W795;
wire W796;
wire W797;
wire W798;
wire W799;
wire W800;
wire W801;
wire W802;
wire W803;
wire W804;
wire W805;
wire W806;
wire W807;
wire W808;
wire W809;
wire W810;
wire W811;
wire W812;
wire W813;
wire W814;
wire W815;
wire W816;
wire W817;
wire W818;
wire W819;
wire W820;
wire W821;
wire W822;
wire W823;
wire W824;
wire W825;
wire W826;
wire W827;
wire W828;
wire W829;
wire W830;
wire W831;
wire W832;
wire W833;
wire W834;
wire W835;
wire W836;
wire W837;
wire W838;
wire W839;
wire W840;
wire W841;
wire W842;
wire W843;
wire W844;
wire W845;
wire W846;
wire W847;
wire W848;
wire W849;
wire W850;
wire W851;
wire W852;
wire W853;
wire W854;
wire W855;
wire W856;
wire W857;
wire W858;
wire W859;
wire W860;
wire W861;
wire W862;
wire W863;
wire W864;
wire W865;
wire W866;
wire W867;
wire W868;
wire W869;
wire W870;
wire W871;
wire W872;
wire W873;
wire W874;
wire W875;
wire W876;
wire W877;
wire W878;
wire W879;
wire W880;
wire W881;
wire W882;
wire W883;
wire W884;
wire W885;
wire W886;
wire W887;
wire W888;
wire W889;
wire W890;
wire W891;
wire W892;
wire W893;
wire W894;
wire W895;
wire W896;
wire W897;
wire W898;
wire W899;
wire W900;
wire W901;
wire W902;
wire W903;
wire W904;
wire W905;
wire W906;
wire W907;
wire W908;
wire W909;
wire W910;
wire W911;
wire W912;
wire W913;
wire W914;
wire W915;
wire W916;
wire W917;
wire W918;
wire W919;
wire W920;
wire W921;
wire W922;
wire W923;
wire W924;
wire W925;
wire W926;
wire W927;
wire W928;
wire W929;
wire W930;
wire W931;
wire W932;
wire W933;
wire W934;
wire W935;
wire W936;
wire W937;
wire W938;
wire W939;
wire W940;
wire W941;
wire W942;
wire W943;
wire W944;
wire W945;
wire W946;
wire W947;
wire W948;
wire W949;
wire W950;
wire W951;
wire W952;
wire W953;
wire W954;
wire W955;
wire W956;
wire W957;
wire W958;
wire W959;
wire W960;
wire W961;
wire W962;
wire W963;
wire W964;
wire W965;
wire W966;
wire W967;
wire W968;
wire W969;
wire W970;
wire W971;
wire W972;
wire W973;
wire W974;
wire W975;
wire W976;
wire W977;
wire W978;
wire W979;
wire W980;
wire W981;
wire W982;
wire W983;
wire W984;
wire W985;
wire W986;
wire W987;
wire W988;
wire W989;
wire W990;
wire W991;
wire W992;
wire W993;
wire W994;
wire W995;
wire W996;
wire W997;
wire W998;
wire W999;
wire W1000;
wire W1001;
wire W1002;
wire W1003;
wire W1004;
wire W1005;
wire W1006;
wire W1007;
wire W1008;
wire W1009;
wire W1010;
wire W1011;
wire W1012;
wire W1013;
wire W1014;
wire W1015;
wire W1016;
wire W1017;
wire W1018;
wire W1019;
wire W1020;
wire W1021;
wire W1022;
wire W1023;
wire W1024;
wire W1025;
wire W1026;
wire W1027;
wire W1028;
wire W1029;
wire W1030;
wire W1031;
wire W1032;
wire W1033;
wire W1034;
wire W1035;
wire W1036;
wire W1037;
wire W1038;
wire W1039;
wire W1040;
wire W1041;
wire W1042;
wire W1043;
wire W1044;
wire W1045;
wire W1046;
wire W1047;
wire W1048;
wire W1049;
wire W1050;
wire W1051;
wire W1052;
wire W1053;
wire W1054;
wire W1055;
wire W1056;
wire W1057;
wire W1058;
wire W1059;
wire W1060;
wire W1061;
wire W1062;
wire W1063;
wire W1064;
wire W1065;
wire W1066;
wire W1067;
wire W1068;
wire W1069;
wire W1070;
wire W1071;
wire W1072;
wire W1073;
wire W1074;
wire W1075;
wire W1076;
wire W1077;
wire W1078;
wire W1079;
wire W1080;
wire W1081;
wire W1082;
wire W1083;
wire W1084;
wire W1085;
wire W1086;
wire W1087;
wire W1088;
wire W1089;
wire W1090;
wire W1091;
wire W1092;
wire W1093;
wire W1094;
wire W1095;
wire W1096;
wire W1097;
wire W1098;
wire W1099;
wire W1100;
wire W1101;
wire W1102;
wire W1103;
wire W1104;
wire W1105;
wire W1106;
wire W1107;
wire W1108;
wire W1109;
wire W1110;
wire W1111;
wire W1112;
wire W1113;
wire W1114;
wire W1115;
wire W1116;
wire W1117;
wire W1118;
wire W1119;
wire W1120;
wire W1121;
wire W1122;
wire W1123;
wire W1124;
wire W1125;
wire W1126;
wire W1127;
wire W1128;
wire W1129;
wire W1130;
wire W1131;
wire W1132;
wire W1133;
wire W1134;
wire W1135;
wire W1136;
wire W1137;
wire W1138;
wire W1139;
wire W1140;
wire W1141;
wire W1142;
wire W1143;
wire W1144;
wire W1145;
wire W1146;
wire W1147;
wire W1148;
wire W1149;
wire W1150;
wire W1151;
wire W1152;
wire W1153;
wire W1154;
wire W1155;
wire W1156;
wire W1157;
wire W1158;
wire W1159;
wire W1160;
wire W1161;
wire W1162;
wire W1163;
wire W1164;
wire W1165;
wire W1166;
wire W1167;
wire W1168;
wire W1169;
wire W1170;
wire W1171;
wire W1172;
wire W1173;
wire W1174;
wire W1175;
wire W1176;
wire W1177;
wire W1178;
wire W1179;
wire W1180;
wire W1181;
wire W1182;
wire W1183;
wire W1184;
wire W1185;
wire W1186;
wire W1187;
wire W1188;
wire W1189;
wire W1190;
wire W1191;
wire W1192;
wire W1193;
wire W1194;
wire W1195;
wire W1196;
wire W1197;
wire W1198;
wire W1199;
wire W1200;
wire W1201;
wire W1202;
wire W1203;
wire W1204;
wire W1205;
wire W1206;
wire W1207;
wire W1208;
wire W1209;
wire W1210;
wire W1211;
wire W1212;
wire W1213;
wire W1214;
wire W1215;
wire W1216;
wire W1217;
wire W1218;
wire W1219;
wire W1220;
wire W1221;
wire W1222;
wire W1223;
wire W1224;
wire W1225;
wire W1226;
wire W1227;
wire W1228;
wire W1229;
wire W1230;
wire W1231;
wire W1232;
wire W1233;
wire W1234;
wire W1235;
wire W1236;
wire W1237;
wire W1238;
wire W1239;
wire W1240;
wire W1241;
wire W1242;
wire W1243;
wire W1244;
wire W1245;
wire W1246;
wire W1247;
wire W1248;
wire W1249;
wire W1250;
wire W1251;
wire W1252;
wire W1253;
wire W1254;
wire W1255;
wire W1256;
wire W1257;
wire W1258;
wire W1259;
wire W1260;
wire W1261;
wire W1262;
wire W1263;
wire W1264;
wire W1265;
wire W1266;
wire W1267;
wire W1268;
wire W1269;
wire W1270;
wire W1271;
wire W1272;
wire W1273;
wire W1274;
wire W1275;
wire W1276;
wire W1277;
wire W1278;
wire W1279;
wire W1280;
wire W1281;
wire W1282;
wire W1283;
wire W1284;
wire W1285;
wire W1286;
wire W1287;
wire W1288;
wire W1289;
wire W1290;
wire W1291;
wire W1292;
wire W1293;
wire W1294;
wire W1295;
wire W1296;
wire W1297;
wire W1298;
wire W1299;
wire W1300;
wire W1301;
wire W1302;
wire W1303;
wire W1304;
wire W1305;
wire W1306;
wire W1307;
wire W1308;
wire W1309;
wire W1310;
wire W1311;
wire W1312;
wire W1313;
wire W1314;
wire W1315;
wire W1316;
wire W1317;
wire W1318;
wire W1319;
wire W1320;
wire W1321;
wire W1322;
wire W1323;
wire W1324;
wire W1325;
wire W1326;
wire W1327;
wire W1328;
wire W1329;
wire W1330;
wire W1331;
wire W1332;
wire W1333;
wire W1334;
wire W1335;
wire W1336;
wire W1337;
wire W1338;
wire W1339;
wire W1340;
wire W1341;
wire W1342;
wire W1343;
wire W1344;
wire W1345;
wire W1346;
wire W1347;
wire W1348;
wire W1349;
wire W1350;
wire W1351;
wire W1352;
wire W1353;
wire W1354;
wire W1355;
wire W1356;
wire W1357;
wire W1358;
wire W1359;
wire W1360;
wire W1361;
wire W1362;
wire W1363;
wire W1364;
wire W1365;
wire W1366;
wire W1367;
wire W1368;
wire W1369;
wire W1370;
wire W1371;
wire W1372;
wire W1373;
wire W1374;
wire W1375;
wire W1376;
wire W1377;
wire W1378;
wire W1379;
wire W1380;
wire W1381;
wire W1382;
wire W1383;
wire W1384;
wire W1385;
wire W1386;
wire W1387;
wire W1388;
wire W1389;
wire W1390;
wire W1391;
wire W1392;
wire W1393;
wire W1394;
wire W1395;
wire W1396;
wire W1397;
wire W1398;
wire W1399;
wire W1400;
wire W1401;
wire W1402;
wire W1403;
wire W1404;
wire W1405;
wire W1406;
wire W1407;
wire W1408;
wire W1409;
wire W1410;
wire W1411;
wire W1412;
wire W1413;
wire W1414;
wire W1415;
wire W1416;
wire W1417;
wire W1418;
wire W1419;
wire W1420;
wire W1421;
wire W1422;
wire W1423;
wire W1424;
wire W1425;
wire W1426;
wire W1427;
wire W1428;
wire W1429;
wire W1430;
wire W1431;
wire W1432;
wire W1433;
wire W1434;
wire W1435;
wire W1436;
wire W1437;
wire W1438;
wire W1439;
wire W1440;
wire W1441;
wire W1442;
wire W1443;
wire W1444;
wire W1445;
wire W1446;
wire W1447;
wire W1448;
wire W1449;
wire W1450;
wire W1451;
wire W1452;
wire W1453;
wire W1454;
wire W1455;
wire W1456;
wire W1457;
wire W1458;
wire W1459;
wire W1460;
wire W1461;
wire W1462;
wire W1463;
wire W1464;
wire W1465;
wire W1466;
wire W1467;
wire W1468;
wire W1469;
wire W1470;
wire W1471;
wire W1472;
wire W1473;
wire W1474;
wire W1475;
wire W1476;
wire W1477;
wire W1478;
wire W1479;
wire W1480;
wire W1481;
wire W1482;
wire W1483;
wire W1484;
wire W1485;
wire W1486;
wire W1487;
wire W1488;
wire W1489;
wire W1490;
wire W1491;
wire W1492;
wire W1493;
wire W1494;
wire W1495;
wire W1496;
wire W1497;
wire W1498;
wire W1499;
wire W1500;
wire W1501;
wire W1502;
wire W1503;
wire W1504;
wire W1505;
wire W1506;
wire W1507;
wire W1508;
wire W1509;
wire W1510;
wire W1511;
wire W1512;
wire W1513;
wire W1514;
wire W1515;
wire W1516;
wire W1517;
wire W1518;
wire W1519;
wire W1520;
wire W1521;
wire W1522;
wire W1523;
wire W1524;
wire W1525;
wire W1526;
wire W1527;
wire W1528;
wire W1529;
wire W1530;
wire W1531;
wire W1532;
wire W1533;
wire W1534;
wire W1535;
wire W1536;
wire W1537;
wire W1538;
wire W1539;
wire W1540;
wire W1541;
wire W1542;
wire W1543;
wire W1544;
wire W1545;
wire W1546;
wire W1547;
wire W1548;
wire W1549;
wire W1550;
wire W1551;
wire W1552;
wire W1553;
wire W1554;
wire W1555;
wire W1556;
wire W1557;
wire W1558;
wire W1559;
wire W1560;
wire W1561;
wire W1562;
wire W1563;
wire W1564;
wire W1565;
wire W1566;
wire W1567;
wire W1568;
wire W1569;
wire W1570;
wire W1571;
wire W1572;
wire W1573;
wire W1574;
wire W1575;
wire W1576;
wire W1577;
wire W1578;
wire W1579;
wire W1580;
wire W1581;
wire W1582;
wire W1583;
wire W1584;
wire W1585;
wire W1586;
wire W1587;
wire W1588;
wire W1589;
wire W1590;
wire W1591;
wire W1592;
wire W1593;
wire W1594;
wire W1595;
wire W1596;
wire W1597;
wire W1598;
wire W1599;
wire W1600;
wire W1601;
wire W1602;
wire W1603;
wire W1604;
wire W1605;
wire W1606;
wire W1607;
wire W1608;
wire W1609;
wire W1610;
wire W1611;
wire W1612;
wire W1613;
wire W1614;
wire W1615;
wire W1616;
wire W1617;
wire W1618;
wire W1619;
wire W1620;
wire W1621;
wire W1622;
wire W1623;
wire W1624;
wire W1625;
wire W1626;
wire W1627;
wire W1628;
wire W1629;
wire W1630;
wire W1631;
wire W1632;
wire W1633;
wire W1634;
wire W1635;
wire W1636;
wire W1637;
wire W1638;
wire W1639;
wire W1640;
wire W1641;
wire W1642;
wire W1643;
wire W1644;
wire W1645;
wire W1646;
wire W1647;
wire W1648;
wire W1649;
wire W1650;
wire W1651;
wire W1652;
wire W1653;
wire W1654;
wire W1655;
wire W1656;
wire W1657;
wire W1658;
wire W1659;
wire W1660;
wire W1661;
wire W1662;
wire W1663;
wire W1664;
wire W1665;
wire W1666;
wire W1667;
wire W1668;
wire W1669;
wire W1670;
wire W1671;
wire W1672;
wire W1673;
wire W1674;
wire W1675;
wire W1676;
wire W1677;
wire W1678;
wire W1679;
wire W1680;
wire W1681;
wire W1682;
wire W1683;
wire W1684;
wire W1685;
wire W1686;
wire W1687;
wire W1688;
wire W1689;
wire W1690;
wire W1691;
wire W1692;
wire W1693;
wire W1694;
wire W1695;
wire W1696;
wire W1697;
wire W1698;
wire W1699;
wire W1700;
wire W1701;
wire W1702;
wire W1703;
wire W1704;
wire W1705;
wire W1706;
wire W1707;
wire W1708;
wire W1709;
wire W1710;
wire W1711;
wire W1712;
wire W1713;
wire W1714;
wire W1715;
wire W1716;
wire W1717;
wire W1718;
wire W1719;
wire W1720;
wire W1721;
wire W1722;
wire W1723;
wire W1724;
wire W1725;
wire W1726;
wire W1727;
wire W1728;
wire W1729;
wire W1730;
wire W1731;
wire W1732;
wire W1733;
wire W1734;
wire W1735;
wire W1736;
wire W1737;
wire W1738;
wire W1739;
wire W1740;
wire W1741;
wire W1742;
wire W1743;
wire W1744;
wire W1745;
wire W1746;
wire W1747;
wire W1748;
wire W1749;
wire W1750;
wire W1751;
wire W1752;
wire W1753;
wire W1754;
wire W1755;
wire W1756;
wire W1757;
wire W1758;
wire W1759;
wire W1760;
wire W1761;
wire W1762;
wire W1763;
wire W1764;
wire W1765;
wire W1766;
wire W1767;
wire W1768;
wire W1769;
wire W1770;
wire W1771;
wire W1772;
wire W1773;
wire W1774;
wire W1775;
wire W1776;
wire W1777;
wire W1778;
wire W1779;
wire W1780;
wire W1781;
wire W1782;
wire W1783;
wire W1784;
wire W1785;
wire W1786;
wire W1787;
wire W1788;
wire W1789;
wire W1790;
wire W1791;
wire W1792;
wire W1793;
wire W1794;
wire W1795;
wire W1796;
wire W1797;
wire W1798;
wire W1799;
wire W1800;
wire W1801;
wire W1802;
wire W1803;
wire W1804;
wire W1805;
wire W1806;
wire W1807;
wire W1808;
wire W1809;
wire W1810;
wire W1811;
wire W1812;
wire W1813;
wire W1814;
wire W1815;
wire W1816;
wire W1817;
wire W1818;
wire W1819;
wire W1820;
wire W1821;
wire W1822;
wire W1823;
wire W1824;
wire W1825;
wire W1826;
wire W1827;
wire W1828;
wire W1829;
wire W1830;
wire W1831;
wire W1832;
wire W1833;
wire W1834;
wire W1835;
wire W1836;
wire W1837;
wire W1838;
wire W1839;
wire W1840;
wire W1841;
wire W1842;
wire W1843;
wire W1844;
wire W1845;
wire W1846;
wire W1847;
wire W1848;
wire W1849;
wire W1850;
wire W1851;
wire W1852;
wire W1853;
wire W1854;
wire W1855;
wire W1856;
wire W1857;
wire W1858;
wire W1859;
wire W1860;
wire W1861;
wire W1862;
wire W1863;
wire W1864;
wire W1865;
wire W1866;
wire W1867;
wire W1868;
wire W1869;
wire W1870;
wire W1871;
wire W1872;
wire W1873;
wire W1874;
wire W1875;
wire W1876;
wire W1877;
wire W1878;
wire W1879;
wire W1880;
wire W1881;
wire W1882;
wire W1883;
wire W1884;
wire W1885;
wire W1886;
wire W1887;
wire W1888;
wire W1889;
wire W1890;
wire W1891;
wire W1892;
wire W1893;
wire W1894;
wire W1895;
wire W1896;
wire W1897;
wire W1898;
wire W1899;
wire W1900;
wire W1901;
wire W1902;
wire W1903;
wire W1904;
wire W1905;
wire W1906;
wire W1907;
wire W1908;
wire W1909;
wire W1910;
wire W1911;
wire W1912;
wire W1913;
wire W1914;
wire W1915;
wire W1916;
wire W1917;
wire W1918;
wire W1919;
wire W1920;
wire W1921;
wire W1922;
wire W1923;
wire W1924;
wire W1925;
wire W1926;
wire W1927;
wire W1928;
wire W1929;
wire W1930;
wire W1931;
wire W1932;
wire W1933;
wire W1934;
wire W1935;
wire W1936;
wire W1937;
wire W1938;
wire W1939;
wire W1940;
wire W1941;
wire W1942;
wire W1943;
wire W1944;
wire W1945;
wire W1946;
wire W1947;
wire W1948;
wire W1949;
wire W1950;
wire W1951;
wire W1952;
wire W1953;
wire W1954;
wire W1955;
wire W1956;
wire W1957;
wire W1958;
wire W1959;
wire W1960;
wire W1961;
wire W1962;
wire W1963;
wire W1964;
wire W1965;
wire W1966;
wire W1967;
wire W1968;
wire W1969;
wire W1970;
wire W1971;
wire W1972;
wire W1973;
wire W1974;
wire W1975;
wire W1976;
wire W1977;
wire W1978;
wire W1979;
wire W1980;
wire W1981;
wire W1982;
wire W1983;
wire W1984;
wire W1985;
wire W1986;
wire W1987;
wire W1988;
wire W1989;
wire W1990;
wire W1991;
wire W1992;
wire W1993;
wire W1994;
wire W1995;
wire W1996;
wire W1997;
wire W1998;
wire W1999;
wire W2000;
wire W2001;
wire W2002;
wire W2003;
wire W2004;
wire W2005;
wire W2006;
wire W2007;
wire W2008;
wire W2009;
wire W2010;
wire W2011;
wire W2012;
wire W2013;
wire W2014;
wire W2015;
wire W2016;
wire W2017;
wire W2018;
wire W2019;
wire W2020;
wire W2021;
wire W2022;
wire W2023;
wire W2024;
wire W2025;
wire W2026;
wire W2027;
wire W2028;
wire W2029;
wire W2030;
wire W2031;
wire W2032;
wire W2033;
wire W2034;
wire W2035;
wire W2036;
wire W2037;
wire W2038;
wire W2039;
wire W2040;
wire W2041;
wire W2042;
wire W2043;
wire W2044;
wire W2045;
wire W2046;
wire W2047;
wire W2048;
wire W2049;
wire W2050;
wire W2051;
wire W2052;
wire W2053;
wire W2054;
wire W2055;
wire W2056;
wire W2057;
wire W2058;
wire W2059;
wire W2060;
wire W2061;
wire W2062;
wire W2063;
wire W2064;
wire W2065;
wire W2066;
wire W2067;
wire W2068;
wire W2069;
wire W2070;
wire W2071;
wire W2072;
wire W2073;
wire W2074;
wire W2075;
wire W2076;
wire W2077;
wire W2078;
wire W2079;
wire W2080;
wire W2081;
wire W2082;
wire W2083;
wire W2084;
wire W2085;
wire W2086;
wire W2087;
wire W2088;
wire W2089;
wire W2090;
wire W2091;
wire W2092;
wire W2093;
wire W2094;
wire W2095;
wire W2096;
wire W2097;
wire W2098;
wire W2099;
wire W2100;
wire W2101;
wire W2102;
wire W2103;
wire W2104;
wire W2105;
wire W2106;
wire W2107;
wire W2108;
wire W2109;
wire W2110;
wire W2111;
wire W2112;
wire W2113;
wire W2114;
wire W2115;
wire W2116;
wire W2117;
wire W2118;
wire W2119;
wire W2120;
wire W2121;
wire W2122;
wire W2123;
wire W2124;
wire W2125;
wire W2126;
wire W2127;
wire W2128;
wire W2129;
wire W2130;
wire W2131;
wire W2132;
wire W2133;
wire W2134;
wire W2135;
wire W2136;
wire W2137;
wire W2138;
wire W2139;
wire W2140;
wire W2141;
wire W2142;
wire W2143;
wire W2144;
wire W2145;
wire W2146;
wire W2147;
wire W2148;
wire W2149;
wire W2150;
wire W2151;
wire W2152;
wire W2153;
wire W2154;
wire W2155;
wire W2156;
wire W2157;
wire W2158;
wire W2159;
wire W2160;
wire W2161;
wire W2162;
wire W2163;
wire W2164;
wire W2165;
wire W2166;
wire W2167;
wire W2168;
wire W2169;
wire W2170;
wire W2171;
wire W2172;
wire W2173;
wire W2174;
wire W2175;
wire W2176;
wire W2177;
wire W2178;
wire W2179;
wire W2180;
wire W2181;
wire W2182;
wire W2183;
wire W2184;
wire W2185;
wire W2186;
wire W2187;
wire W2188;
wire W2189;
wire W2190;
wire W2191;
wire W2192;
wire W2193;
wire W2194;
wire W2195;
wire W2196;
wire W2197;
wire W2198;
wire W2199;
wire W2200;
wire W2201;
wire W2202;
wire W2203;
wire W2204;
wire W2205;
wire W2206;
wire W2207;
wire W2208;
wire W2209;
wire W2210;
wire W2211;
wire W2212;
wire W2213;
wire W2214;
wire W2215;
wire W2216;
wire W2217;
wire W2218;
wire W2219;
wire W2220;
wire W2221;
wire W2222;
wire W2223;
wire W2224;
wire W2225;
wire W2226;
wire W2227;
wire W2228;
wire W2229;
wire W2230;
wire W2231;
wire W2232;
wire W2233;
wire W2234;
wire W2235;
wire W2236;
wire W2237;
wire W2238;
wire W2239;
wire W2240;
wire W2241;
wire W2242;
wire W2243;
wire W2244;
wire W2245;
wire W2246;
wire W2247;
wire W2248;
wire W2249;
wire W2250;
wire W2251;
wire W2252;
wire W2253;
wire W2254;
wire W2255;
wire W2256;
wire W2257;
wire W2258;
wire W2259;
wire W2260;
wire W2261;
wire W2262;
wire W2263;
wire W2264;
wire W2265;
wire W2266;
wire W2267;
wire W2268;
wire W2269;
wire W2270;
wire W2271;
wire W2272;
wire W2273;
wire W2274;
wire W2275;
wire W2276;
wire W2277;
wire W2278;
wire W2279;
wire W2280;
wire W2281;
wire W2282;
wire W2283;
wire W2284;
wire W2285;
wire W2286;
wire W2287;
wire W2288;
wire W2289;
wire W2290;
wire W2291;
wire W2292;
wire W2293;
wire W2294;
wire W2295;
wire W2296;
wire W2297;
wire W2298;
wire W2299;
wire W2300;
wire W2301;
wire W2302;
wire W2303;
wire W2304;
wire W2305;
wire W2306;
wire W2307;
wire W2308;
wire W2309;
wire W2310;
wire W2311;
wire W2312;
wire W2313;
wire W2314;
wire W2315;
wire W2316;
wire W2317;
wire W2318;
wire W2319;
wire W2320;
wire W2321;
wire W2322;
wire W2323;
wire W2324;
wire W2325;
wire W2326;
wire W2327;
wire W2328;
wire W2329;
wire W2330;
wire W2331;
wire W2332;
wire W2333;
wire W2334;
wire W2335;
wire W2336;
wire W2337;
wire W2338;
wire W2339;
wire W2340;
wire W2341;
wire W2342;
wire W2343;
wire W2344;
wire W2345;
wire W2346;
wire W2347;
wire W2348;
wire W2349;
wire W2350;
wire W2351;
wire W2352;
wire W2353;
wire W2354;
wire W2355;
wire W2356;
wire W2357;
wire W2358;
wire W2359;
wire W2360;
wire W2361;
wire W2362;
wire W2363;
wire W2364;
wire W2365;
wire W2366;
wire W2367;
wire W2368;
wire W2369;
wire W2370;
wire W2371;
wire W2372;
wire W2373;
wire W2374;
wire W2375;
wire W2376;
wire W2377;
wire W2378;
wire W2379;
wire W2380;
wire W2381;
wire W2382;
wire W2383;
wire W2384;
wire W2385;
wire W2386;
wire W2387;
wire W2388;
wire W2389;
wire W2390;
wire W2391;
wire W2392;
wire W2393;
wire W2394;
wire W2395;
wire W2396;
wire W2397;
wire W2398;
wire W2399;
wire W2400;
wire W2401;
wire W2402;
wire W2403;
wire W2404;
wire W2405;
wire W2406;
wire W2407;
wire W2408;
wire W2409;
wire W2410;
wire W2411;
wire W2412;
wire W2413;
wire W2414;
wire W2415;
wire W2416;
wire W2417;
wire W2418;
wire W2419;
wire W2420;
wire W2421;
wire W2422;
wire W2423;
wire W2424;
wire W2425;
wire W2426;
wire W2427;
wire W2428;
wire W2429;
wire W2430;
wire W2431;
wire W2432;
wire W2433;
wire W2434;
wire W2435;
wire W2436;
wire W2437;
wire W2438;
wire W2439;
wire W2440;
wire W2441;
wire W2442;
wire W2443;
wire W2444;
wire W2445;
wire W2446;
wire W2447;
wire W2448;
wire W2449;
wire W2450;
wire W2451;
wire W2452;
wire W2453;
wire W2454;
wire W2455;
wire W2456;
wire W2457;
wire W2458;
wire W2459;
wire W2460;
wire W2461;
wire W2462;
wire W2463;
wire W2464;
wire W2465;
wire W2466;
wire W2467;
wire W2468;
wire W2469;
wire W2470;
wire W2471;
wire W2472;
wire W2473;
wire W2474;
wire W2475;
wire W2476;
wire W2477;
wire W2478;
wire W2479;
wire W2480;
wire W2481;
wire W2482;
wire W2483;
wire W2484;
wire W2485;
wire W2486;
wire W2487;
wire W2488;
wire W2489;
wire W2490;
wire W2491;
wire W2492;
wire W2493;
wire W2494;
wire W2495;
wire W2496;
wire W2497;
wire W2498;
wire W2499;
wire W2500;
wire W2501;
wire W2502;
wire W2503;
wire W2504;
wire W2505;
wire W2506;
wire W2507;
wire W2508;
wire W2509;
wire W2510;
wire W2511;
wire W2512;
wire W2513;
wire W2514;
wire W2515;
wire W2516;
wire W2517;
wire W2518;
wire W2519;
wire W2520;
wire W2521;
wire W2522;
wire W2523;
wire W2524;
wire W2525;
wire W2526;
wire W2527;
wire W2528;
wire W2529;
wire W2530;
wire W2531;
wire W2532;
wire W2533;
wire W2534;
wire W2535;
wire W2536;
wire W2537;
wire W2538;
wire W2539;
wire W2540;
wire W2541;
wire W2542;
wire W2543;
wire W2544;
wire W2545;
wire W2546;
wire W2547;
wire W2548;
wire W2549;
wire W2550;
wire W2551;
wire W2552;
wire W2553;
wire W2554;
wire W2555;
wire W2556;
wire W2557;
wire W2558;
wire W2559;
wire W2560;
wire W2561;
wire W2562;
wire W2563;
wire W2564;
wire W2565;
wire W2566;
wire W2567;
wire W2568;
wire W2569;
wire W2570;
wire W2571;
wire W2572;
wire W2573;
wire W2574;
wire W2575;
wire W2576;
wire W2577;
wire W2578;
wire W2579;
wire W2580;
wire W2581;
wire W2582;
wire W2583;
wire W2584;
wire W2585;
wire W2586;
wire W2587;
wire W2588;
wire W2589;
wire W2590;
wire W2591;
wire W2592;
wire W2593;
wire W2594;
wire W2595;
wire W2596;
wire W2597;
wire W2598;
wire W2599;
wire W2600;
wire W2601;
wire W2602;
wire W2603;
wire W2604;
wire W2605;
wire W2606;
wire W2607;
wire W2608;
wire W2609;
wire W2610;
wire W2611;
wire W2612;
wire W2613;
wire W2614;
wire W2615;
wire W2616;
wire W2617;
wire W2618;
wire W2619;
wire W2620;
wire W2621;
wire W2622;
wire W2623;
wire W2624;
wire W2625;
wire W2626;
wire W2627;
wire W2628;
wire W2629;
wire W2630;
wire W2631;
wire W2632;
wire W2633;
wire W2634;
wire W2635;
wire W2636;
wire W2637;
wire W2638;
wire W2639;
wire W2640;
wire W2641;
wire W2642;
wire W2643;
wire W2644;
wire W2645;
wire W2646;
wire W2647;
wire W2648;
wire W2649;
wire W2650;
wire W2651;
wire W2652;
wire W2653;
wire W2654;
wire W2655;
wire W2656;
wire W2657;
wire W2658;
wire W2659;
wire W2660;
wire W2661;
wire W2662;
wire W2663;
wire W2664;
wire W2665;
wire W2666;
wire W2667;
wire W2668;
wire W2669;
wire W2670;
wire W2671;
wire W2672;
wire W2673;
wire W2674;
wire W2675;
wire W2676;
wire W2677;
wire W2678;
wire W2679;
wire W2680;
wire W2681;
wire W2682;
wire W2683;
wire W2684;
wire W2685;
wire W2686;
wire W2687;
wire W2688;
wire W2689;
wire W2690;
wire W2691;
wire W2692;
wire W2693;
wire W2694;
wire W2695;
wire W2696;
wire W2697;
wire W2698;
wire W2699;
wire W2700;
wire W2701;
wire W2702;
wire W2703;
wire W2704;
wire W2705;
wire W2706;
wire W2707;
wire W2708;
wire W2709;
wire W2710;
wire W2711;
wire W2712;
wire W2713;
wire W2714;
wire W2715;
wire W2716;
wire W2717;
wire W2718;
wire W2719;
wire W2720;
wire W2721;
wire W2722;
wire W2723;
wire W2724;
wire W2725;
wire W2726;
wire W2727;
wire W2728;
wire W2729;
wire W2730;
wire W2731;
wire W2732;
wire W2733;
wire W2734;
wire W2735;
wire W2736;
wire W2737;
wire W2738;
wire W2739;
wire W2740;
wire W2741;
wire W2742;
wire W2743;
wire W2744;
wire W2745;
wire W2746;
wire W2747;
wire W2748;
wire W2749;
wire W2750;
wire W2751;
wire W2752;
wire W2753;
wire W2754;
wire W2755;
wire W2756;
wire W2757;
wire W2758;
wire W2759;
wire W2760;
wire W2761;
wire W2762;
wire W2763;
wire W2764;
wire W2765;
wire W2766;
wire W2767;
wire W2768;
wire W2769;
wire W2770;
wire W2771;
wire W2772;
wire W2773;
wire W2774;
wire W2775;
wire W2776;
wire W2777;
wire W2778;
wire W2779;
wire W2780;
wire W2781;
wire W2782;
wire W2783;
wire W2784;
wire W2785;
wire W2786;
wire W2787;
wire W2788;
wire W2789;
wire W2790;
wire W2791;
wire W2792;
wire W2793;
wire W2794;
wire W2795;
wire W2796;
wire W2797;
wire W2798;
wire W2799;
wire W2800;
wire W2801;
wire W2802;
wire W2803;
wire W2804;
wire W2805;
wire W2806;
wire W2807;
wire W2808;
wire W2809;
wire W2810;
wire W2811;
wire W2812;
wire W2813;
wire W2814;
wire W2815;
wire W2816;
wire W2817;
wire W2818;
wire W2819;
wire W2820;
wire W2821;
wire W2822;
wire W2823;
wire W2824;
wire W2825;
wire W2826;
wire W2827;
wire W2828;
wire W2829;
wire W2830;
wire W2831;
wire W2832;
wire W2833;
wire W2834;
wire W2835;
wire W2836;
wire W2837;
wire W2838;
wire W2839;
wire W2840;
wire W2841;
wire W2842;
wire W2843;
wire W2844;
wire W2845;
wire W2846;
wire W2847;
wire W2848;
wire W2849;
wire W2850;
wire W2851;
wire W2852;
wire W2853;
wire W2854;
wire W2855;
wire W2856;
wire W2857;
wire W2858;
wire W2859;
wire W2860;
wire W2861;
wire W2862;
wire W2863;
wire W2864;
wire W2865;
wire W2866;
wire W2867;
wire W2868;
wire W2869;
wire W2870;
wire W2871;
wire W2872;
wire W2873;
wire W2874;
wire W2875;
wire W2876;
wire W2877;
wire W2878;
wire W2879;
wire W2880;
wire W2881;
wire W2882;
wire W2883;
wire W2884;
wire W2885;
wire W2886;
wire W2887;
wire W2888;
wire W2889;
wire W2890;
wire W2891;
wire W2892;
wire W2893;
wire W2894;
wire W2895;
wire W2896;
wire W2897;
wire W2898;
wire W2899;
wire W2900;
wire W2901;
wire W2902;
wire W2903;
wire W2904;
wire W2905;
wire W2906;
wire W2907;
wire W2908;
wire W2909;
wire W2910;
wire W2911;
wire W2912;
wire W2913;
wire W2914;
wire W2915;
wire W2916;
wire W2917;
wire W2918;
wire W2919;
wire W2920;
wire W2921;
wire W2922;
wire W2923;
wire W2924;
wire W2925;
wire W2926;
wire W2927;
wire W2928;
wire W2929;
wire W2930;
wire W2931;
wire W2932;
wire W2933;
wire W2934;
wire W2935;
wire W2936;
wire W2937;
wire W2938;
wire W2939;
wire W2940;
wire W2941;
wire W2942;
wire W2943;
wire W2944;
wire W2945;
wire W2946;
wire W2947;
wire W2948;
wire W2949;
wire W2950;
wire W2951;
wire W2952;
wire W2953;
wire W2954;
wire W2955;
wire W2956;
wire W2957;
wire W2958;
wire W2959;
wire W2960;
wire W2961;
wire W2962;
wire W2963;
wire W2964;
wire W2965;
wire W2966;
wire W2967;
wire W2968;
wire W2969;
wire W2970;
wire W2971;
wire W2972;
wire W2973;
wire W2974;
wire W2975;
wire W2976;
wire W2977;
wire W2978;
wire W2979;
wire W2980;
wire W2981;
wire W2982;
wire W2983;
wire W2984;
wire W2985;
wire W2986;
wire W2987;
wire W2988;
wire W2989;
wire W2990;
wire W2991;
wire W2992;
wire W2993;
wire W2994;
wire W2995;
wire W2996;
wire W2997;
wire W2998;
wire W2999;
wire W3000;
wire W3001;
wire W3002;
wire W3003;
wire W3004;
wire W3005;
wire W3006;
wire W3007;
wire W3008;
wire W3009;
wire W3010;
wire W3011;
wire W3012;
wire W3013;
wire W3014;
wire W3015;
wire W3016;
wire W3017;
wire W3018;
wire W3019;
wire W3020;
wire W3021;
wire W3022;
wire W3023;
wire W3024;
wire W3025;
wire W3026;
wire W3027;
wire W3028;
wire W3029;
wire W3030;
wire W3031;
wire W3032;
wire W3033;
wire W3034;
wire W3035;
wire W3036;
wire W3037;
wire W3038;
wire W3039;
wire W3040;
wire W3041;
wire W3042;
wire W3043;
wire W3044;
wire W3045;
wire W3046;
wire W3047;
wire W3048;
wire W3049;
wire W3050;
wire W3051;
wire W3052;
wire W3053;
wire W3054;
wire W3055;
wire W3056;
wire W3057;
wire W3058;
wire W3059;
wire W3060;
wire W3061;
wire W3062;
wire W3063;
wire W3064;
wire W3065;
wire W3066;
wire W3067;
wire W3068;
wire W3069;
wire W3070;
wire W3071;
wire W3072;
wire W3073;
wire W3074;
wire W3075;
wire W3076;
wire W3077;
wire W3078;
wire W3079;
wire W3080;
wire W3081;
wire W3082;
wire W3083;
wire W3084;
wire W3085;
wire W3086;
wire W3087;
wire W3088;
wire W3089;
wire W3090;
wire W3091;
wire W3092;
wire W3093;
wire W3094;
wire W3095;
wire W3096;
wire W3097;
wire W3098;
wire W3099;
wire W3100;
wire W3101;
wire W3102;
wire W3103;
wire W3104;
wire W3105;
wire W3106;
wire W3107;
wire W3108;
wire W3109;
wire W3110;
wire W3111;
wire W3112;
wire W3113;
wire W3114;
wire W3115;
wire W3116;
wire W3117;
wire W3118;
wire W3119;
wire W3120;
wire W3121;
wire W3122;
wire W3123;
wire W3124;
wire W3125;
wire W3126;
wire W3127;
wire W3128;
wire W3129;
wire W3130;
wire W3131;
wire W3132;
wire W3133;
wire W3134;
wire W3135;
wire W3136;
wire W3137;
wire W3138;
wire W3139;
wire W3140;
wire W3141;
wire W3142;
wire W3143;
wire W3144;
wire W3145;
wire W3146;
wire W3147;
wire W3148;
wire W3149;
wire W3150;
wire W3151;
wire W3152;
wire W3153;
wire W3154;
wire W3155;
wire W3156;
wire W3157;
wire W3158;
wire W3159;
wire W3160;
wire W3161;
wire W3162;
wire W3163;
wire W3164;
wire W3165;
wire W3166;
wire W3167;
wire W3168;
wire W3169;
wire W3170;
wire W3171;
wire W3172;
wire W3173;
wire W3174;
wire W3175;
wire W3176;
wire W3177;
wire W3178;
wire W3179;
wire W3180;
wire W3181;
wire W3182;
wire W3183;
wire W3184;
wire W3185;
wire W3186;
wire W3187;
wire W3188;
wire W3189;
wire W3190;
wire W3191;
wire W3192;
wire W3193;
wire W3194;
wire W3195;
wire W3196;
wire W3197;
wire W3198;
wire W3199;
wire W3200;
wire W3201;
wire W3202;
wire W3203;
wire W3204;
wire W3205;
wire W3206;
wire W3207;
wire W3208;
wire W3209;
wire W3210;
wire W3211;
wire W3212;
wire W3213;
wire W3214;
wire W3215;
wire W3216;
wire W3217;
wire W3218;
wire W3219;
wire W3220;
wire W3221;
wire W3222;
wire W3223;
wire W3224;
wire W3225;
wire W3226;
wire W3227;
wire W3228;
wire W3229;
wire W3230;
wire W3231;
wire W3232;
wire W3233;
wire W3234;
wire W3235;
wire W3236;
wire W3237;
wire W3238;
wire W3239;
wire W3240;
wire W3241;
wire W3242;
wire W3243;
wire W3244;
wire W3245;
wire W3246;
wire W3247;
wire W3248;
wire W3249;
wire W3250;
wire W3251;
wire W3252;
wire W3253;
wire W3254;
wire W3255;
wire W3256;
wire W3257;
wire W3258;
wire W3259;
wire W3260;
wire W3261;
wire W3262;
wire W3263;
wire W3264;
wire W3265;
wire W3266;
wire W3267;
wire W3268;
wire W3269;
wire W3270;
wire W3271;
wire W3272;
wire W3273;
wire W3274;
wire W3275;
wire W3276;
wire W3277;
wire W3278;
wire W3279;
wire W3280;
wire W3281;
wire W3282;
wire W3283;
wire W3284;
wire W3285;
wire W3286;
wire W3287;
wire W3288;
wire W3289;
wire W3290;
wire W3291;
wire W3292;
wire W3293;
wire W3294;
wire W3295;
wire W3296;
wire W3297;
wire W3298;
wire W3299;
wire W3300;
wire W3301;
wire W3302;
wire W3303;
wire W3304;
wire W3305;
wire W3306;
wire W3307;
wire W3308;
wire W3309;
wire W3310;
wire W3311;
wire W3312;
wire W3313;
wire W3314;
wire W3315;
wire W3316;
wire W3317;
wire W3318;
wire W3319;
wire W3320;
wire W3321;
wire W3322;
wire W3323;
wire W3324;
wire W3325;
wire W3326;
wire W3327;
wire W3328;
wire W3329;
wire W3330;
wire W3331;
wire W3332;
wire W3333;
wire W3334;
wire W3335;
wire W3336;
wire W3337;
wire W3338;
wire W3339;
wire W3340;
wire W3341;
wire W3342;
wire W3343;
wire W3344;
wire W3345;
wire W3346;
wire W3347;
wire W3348;
wire W3349;
wire W3350;
wire W3351;
wire W3352;
wire W3353;
wire W3354;
wire W3355;
wire W3356;
wire W3357;
wire W3358;
wire W3359;
wire W3360;
wire W3361;
wire W3362;
wire W3363;
wire W3364;
wire W3365;
wire W3366;
wire W3367;
wire W3368;
wire W3369;
wire W3370;
wire W3371;
wire W3372;
wire W3373;
wire W3374;
wire W3375;
wire W3376;
wire W3377;
wire W3378;
wire W3379;
wire W3380;
wire W3381;
wire W3382;
wire W3383;
wire W3384;
wire W3385;
wire W3386;
wire W3387;
wire W3388;
wire W3389;
wire W3390;
wire W3391;
wire W3392;
wire W3393;
wire W3394;
wire W3395;
wire W3396;
wire W3397;
wire W3398;
wire W3399;
wire W3400;
wire W3401;
wire W3402;
wire W3403;
wire W3404;
wire W3405;
wire W3406;
wire W3407;
wire W3408;
wire W3409;
wire W3410;
wire W3411;
wire W3412;
wire W3413;
wire W3414;
wire W3415;
wire W3416;
wire W3417;
wire W3418;
wire W3419;
wire W3420;
wire W3421;
wire W3422;
wire W3423;
wire W3424;
wire W3425;
wire W3426;
wire W3427;
wire W3428;
wire W3429;
wire W3430;
wire W3431;
wire W3432;
wire W3433;
wire W3434;
wire W3435;
wire W3436;
wire W3437;
wire W3438;
wire W3439;
wire W3440;
wire W3441;
wire W3442;
wire W3443;
wire W3444;
wire W3445;
wire W3446;
wire W3447;
wire W3448;
wire W3449;
wire W3450;
wire W3451;
wire W3452;
wire W3453;
wire W3454;
wire W3455;
wire W3456;
wire W3457;
wire W3458;
wire W3459;
wire W3460;
wire W3461;
wire W3462;
wire W3463;
wire W3464;
wire W3465;
wire W3466;
wire W3467;
wire W3468;
wire W3469;
wire W3470;
wire W3471;
wire W3472;
wire W3473;
wire W3474;
wire W3475;
wire W3476;
wire W3477;
wire W3478;
wire W3479;
wire W3480;
wire W3481;
wire W3482;
wire W3483;
wire W3484;
wire W3485;
wire W3486;
wire W3487;
wire W3488;
wire W3489;
wire W3490;
wire W3491;
wire W3492;
wire W3493;
wire W3494;
wire W3495;
wire W3496;
wire W3497;
wire W3498;
wire W3499;
wire W3500;
wire W3501;
wire W3502;
wire W3503;
wire W3504;
wire W3505;
wire W3506;
wire W3507;
wire W3508;
wire W3509;
wire W3510;
wire W3511;
wire W3512;
wire W3513;
wire W3514;
wire W3515;
wire W3516;
wire W3517;
wire W3518;
wire W3519;
wire W3520;
wire W3521;
wire W3522;
wire W3523;
wire W3524;
wire W3525;
wire W3526;
wire W3527;
wire W3528;
wire W3529;
wire W3530;
wire W3531;
wire W3532;
wire W3533;
wire W3534;
wire W3535;
wire W3536;
wire W3537;
wire W3538;
wire W3539;
wire W3540;
wire W3541;
wire W3542;
wire W3543;
wire W3544;
wire W3545;
wire W3546;
wire W3547;
wire W3548;
wire W3549;
wire W3550;
wire W3551;
wire W3552;
wire W3553;
wire W3554;
wire W3555;
wire W3556;
wire W3557;
wire W3558;
wire W3559;
wire W3560;
wire W3561;
wire W3562;
wire W3563;
wire W3564;
wire W3565;
wire W3566;
wire W3567;
wire W3568;
wire W3569;
wire W3570;
wire W3571;
wire W3572;
wire W3573;
wire W3574;
wire W3575;
wire W3576;
wire W3577;
wire W3578;
wire W3579;
wire W3580;
wire W3581;
wire W3582;
wire W3583;
wire W3584;
wire W3585;
wire W3586;
wire W3587;
wire W3588;
wire W3589;
wire W3590;
wire W3591;
wire W3592;
wire W3593;
wire W3594;
wire W3595;
wire W3596;
wire W3597;
wire W3598;
wire W3599;
wire W3600;
wire W3601;
wire W3602;
wire W3603;
wire W3604;
wire W3605;
wire W3606;
wire W3607;
wire W3608;
wire W3609;
wire W3610;
wire W3611;
wire W3612;
wire W3613;
wire W3614;
wire W3615;
wire W3616;
wire W3617;
wire W3618;
wire W3619;
wire W3620;
wire W3621;
wire W3622;
wire W3623;
wire W3624;
wire W3625;
wire W3626;
wire W3627;
wire W3628;
wire W3629;
wire W3630;
wire W3631;
wire W3632;
wire W3633;
wire W3634;
wire W3635;
wire W3636;
wire W3637;
wire W3638;
wire W3639;
wire W3640;
wire W3641;
wire W3642;
wire W3643;
wire W3644;
wire W3645;
wire W3646;
wire W3647;
wire W3648;
wire W3649;
wire W3650;
wire W3651;
wire W3652;
wire W3653;
wire W3654;
wire W3655;
wire W3656;
wire W3657;
wire W3658;
wire W3659;
wire W3660;
wire W3661;
wire W3662;
wire W3663;
wire W3664;
wire W3665;
wire W3666;
wire W3667;
wire W3668;
wire W3669;
wire W3670;
wire W3671;
wire W3672;
wire W3673;
wire W3674;
wire W3675;
wire W3676;
wire W3677;
wire W3678;
wire W3679;
wire W3680;
wire W3681;
wire W3682;
wire W3683;
wire W3684;
wire W3685;
wire W3686;
wire W3687;
wire W3688;
wire W3689;
wire W3690;
wire W3691;
wire W3692;
wire W3693;
wire W3694;
wire W3695;
wire W3696;
wire W3697;
wire W3698;
wire W3699;
wire W3700;
wire W3701;
wire W3702;
wire W3703;
wire W3704;
wire W3705;
wire W3706;
wire W3707;
wire W3708;
wire W3709;
wire W3710;
wire W3711;
wire W3712;
wire W3713;
wire W3714;
wire W3715;
wire W3716;
wire W3717;
wire W3718;
wire W3719;
wire W3720;
wire W3721;
wire W3722;
wire W3723;
wire W3724;
wire W3725;
wire W3726;
wire W3727;
wire W3728;
wire W3729;
wire W3730;
wire W3731;
wire W3732;
wire W3733;
wire W3734;
wire W3735;
wire W3736;
wire W3737;
wire W3738;
wire W3739;
wire W3740;
wire W3741;
wire W3742;
wire W3743;
wire W3744;
wire W3745;
wire W3746;
wire W3747;
wire W3748;
wire W3749;
wire W3750;
wire W3751;
wire W3752;
wire W3753;
wire W3754;
wire W3755;
wire W3756;
wire W3757;
wire W3758;
wire W3759;
wire W3760;
wire W3761;
wire W3762;
wire W3763;
wire W3764;
wire W3765;
wire W3766;
wire W3767;
wire W3768;
wire W3769;
wire W3770;
wire W3771;
wire W3772;
wire W3773;
wire W3774;
wire W3775;
wire W3776;
wire W3777;
wire W3778;
wire W3779;
wire W3780;
wire W3781;
wire W3782;
wire W3783;
wire W3784;
wire W3785;
wire W3786;
wire W3787;
wire W3788;
wire W3789;
wire W3790;
wire W3791;
wire W3792;
wire W3793;
wire W3794;
wire W3795;
wire W3796;
wire W3797;
wire W3798;
wire W3799;
wire W3800;
wire W3801;
wire W3802;
wire W3803;
wire W3804;
wire W3805;
wire W3806;
wire W3807;
wire W3808;
wire W3809;
wire W3810;
wire W3811;
wire W3812;
wire W3813;
wire W3814;
wire W3815;
wire W3816;
wire W3817;
wire W3818;
wire W3819;
wire W3820;
wire W3821;
wire W3822;
wire W3823;
wire W3824;
wire W3825;
wire W3826;
wire W3827;
wire W3828;
wire W3829;
wire W3830;
wire W3831;
wire W3832;
wire W3833;
wire W3834;
wire W3835;
wire W3836;
wire W3837;
wire W3838;
wire W3839;
wire W3840;
wire W3841;
wire W3842;
wire W3843;
wire W3844;
wire W3845;
wire W3846;
wire W3847;
wire W3848;
wire W3849;
wire W3850;
wire W3851;
wire W3852;
wire W3853;
wire W3854;
wire W3855;
wire W3856;
wire W3857;
wire W3858;
wire W3859;
wire W3860;
wire W3861;
wire W3862;
wire W3863;
wire W3864;
wire W3865;
wire W3866;
wire W3867;
wire W3868;
wire W3869;
wire W3870;
wire W3871;
wire W3872;
wire W3873;
wire W3874;
wire W3875;
wire W3876;
wire W3877;
wire W3878;
wire W3879;
wire W3880;
wire W3881;
wire W3882;
wire W3883;
wire W3884;
wire W3885;
wire W3886;
wire W3887;
wire W3888;
wire W3889;
wire W3890;
wire W3891;
wire W3892;
wire W3893;
wire W3894;
wire W3895;
wire W3896;
wire W3897;
wire W3898;
wire W3899;
wire W3900;
wire W3901;
wire W3902;
wire W3903;
wire W3904;
wire W3905;
wire W3906;
wire W3907;
wire W3908;
wire W3909;
wire W3910;
wire W3911;
wire W3912;
wire W3913;
wire W3914;
wire W3915;
wire W3916;
wire W3917;
wire W3918;
wire W3919;
wire W3920;
wire W3921;
wire W3922;
wire W3923;
wire W3924;
wire W3925;
wire W3926;
wire W3927;
wire W3928;
wire W3929;
wire W3930;
wire W3931;
wire W3932;
wire W3933;
wire W3934;
wire W3935;
wire W3936;
wire W3937;
wire W3938;
wire W3939;
wire W3940;
wire W3941;
wire W3942;
wire W3943;
wire W3944;
wire W3945;
wire W3946;
wire W3947;
wire W3948;
wire W3949;
wire W3950;
wire W3951;
wire W3952;
wire W3953;
wire W3954;
wire W3955;
wire W3956;
wire W3957;
wire W3958;
wire W3959;
wire W3960;
wire W3961;
wire W3962;
wire W3963;
wire W3964;
wire W3965;
wire W3966;
wire W3967;
wire W3968;
wire W3969;
wire W3970;
wire W3971;
wire W3972;
wire W3973;
wire W3974;
wire W3975;
wire W3976;
wire W3977;
wire W3978;
wire W3979;
wire W3980;
wire W3981;
wire W3982;
wire W3983;
wire W3984;
wire W3985;
wire W3986;
wire W3987;
wire W3988;
wire W3989;
wire W3990;
wire W3991;
wire W3992;
wire W3993;
wire W3994;
wire W3995;
wire W3996;
wire W3997;
wire W3998;
wire W3999;
wire W4000;
wire W4001;
wire W4002;
wire W4003;
wire W4004;
wire W4005;
wire W4006;
wire W4007;
wire W4008;
wire W4009;
wire W4010;
wire W4011;
wire W4012;
wire W4013;
wire W4014;
wire W4015;
wire W4016;
wire W4017;
wire W4018;
wire W4019;
wire W4020;
wire W4021;
wire W4022;
wire W4023;
wire W4024;
wire W4025;
wire W4026;
wire W4027;
wire W4028;
wire W4029;
wire W4030;
wire W4031;
wire W4032;
wire W4033;
wire W4034;
wire W4035;
wire W4036;
wire W4037;
wire W4038;
wire W4039;
wire W4040;
wire W4041;
wire W4042;
wire W4043;
wire W4044;
wire W4045;
wire W4046;
wire W4047;
wire W4048;
wire W4049;
wire W4050;
wire W4051;
wire W4052;
wire W4053;
wire W4054;
wire W4055;
wire W4056;
wire W4057;
wire W4058;
wire W4059;
wire W4060;
wire W4061;
wire W4062;
wire W4063;
wire W4064;
wire W4065;
wire W4066;
wire W4067;
wire W4068;
wire W4069;
wire W4070;
wire W4071;
wire W4072;
wire W4073;
wire W4074;
wire W4075;
wire W4076;
wire W4077;
wire W4078;
wire W4079;
wire W4080;
wire W4081;
wire W4082;
wire W4083;
wire W4084;
wire W4085;
wire W4086;
wire W4087;
wire W4088;
wire W4089;
wire W4090;
wire W4091;
wire W4092;
wire W4093;
wire W4094;
wire W4095;
wire W4096;
wire W4097;
wire W4098;
wire W4099;
wire W4100;
wire W4101;
wire W4102;
wire W4103;
wire W4104;
wire W4105;
wire W4106;
wire W4107;
wire W4108;
wire W4109;
wire W4110;
wire W4111;
wire W4112;
wire W4113;
wire W4114;
wire W4115;
wire W4116;
wire W4117;
wire W4118;
wire W4119;
wire W4120;
wire W4121;
wire W4122;
wire W4123;
wire W4124;
wire W4125;
wire W4126;
wire W4127;
wire W4128;
wire W4129;
wire W4130;
wire W4131;
wire W4132;
wire W4133;
wire W4134;
wire W4135;
wire W4136;
wire W4137;
wire W4138;
wire W4139;
wire W4140;
wire W4141;
wire W4142;
wire W4143;
wire W4144;
wire W4145;
wire W4146;
wire W4147;
wire W4148;
wire W4149;
wire W4150;
wire W4151;
wire W4152;
wire W4153;
wire W4154;
wire W4155;
wire W4156;
wire W4157;
wire W4158;
wire W4159;
wire W4160;
wire W4161;
wire W4162;
wire W4163;
wire W4164;
wire W4165;
wire W4166;
wire W4167;
wire W4168;
wire W4169;
wire W4170;
wire W4171;
wire W4172;
wire W4173;
wire W4174;
wire W4175;
wire W4176;
wire W4177;
wire W4178;
wire W4179;
wire W4180;
wire W4181;
wire W4182;
wire W4183;
wire W4184;
wire W4185;
wire W4186;
wire W4187;
wire W4188;
wire W4189;
wire W4190;
wire W4191;
wire W4192;
wire W4193;
wire W4194;
wire W4195;
wire W4196;
wire W4197;
wire W4198;
wire W4199;
wire W4200;
wire W4201;
wire W4202;
wire W4203;
wire W4204;
wire W4205;
wire W4206;
wire W4207;
wire W4208;
wire W4209;
wire W4210;
wire W4211;
wire W4212;
wire W4213;
wire W4214;
wire W4215;
wire W4216;
wire W4217;
wire W4218;
wire W4219;
wire W4220;
wire W4221;
wire W4222;
wire W4223;
wire W4224;
wire W4225;
wire W4226;
wire W4227;
wire W4228;
wire W4229;
wire W4230;
wire W4231;
wire W4232;
wire W4233;
wire W4234;
wire W4235;
wire W4236;
wire W4237;
wire W4238;
wire W4239;
wire W4240;
wire W4241;
wire W4242;
wire W4243;
wire W4244;
wire W4245;
wire W4246;
wire W4247;
wire W4248;
wire W4249;
wire W4250;
wire W4251;
wire W4252;
wire W4253;
wire W4254;
wire W4255;
wire W4256;
wire W4257;
wire W4258;
wire W4259;
wire W4260;
wire W4261;
wire W4262;
wire W4263;
wire W4264;
wire W4265;
wire W4266;
wire W4267;
wire W4268;
wire W4269;
wire W4270;
wire W4271;
wire W4272;
wire W4273;
wire W4274;
wire W4275;
wire W4276;
wire W4277;
wire W4278;
wire W4279;
wire W4280;
wire W4281;
wire W4282;
wire W4283;
wire W4284;
wire W4285;
wire W4286;
wire W4287;
wire W4288;
wire W4289;
wire W4290;
wire W4291;
wire W4292;
wire W4293;
wire W4294;
wire W4295;
wire W4296;
wire W4297;
wire W4298;
wire W4299;
wire W4300;
wire W4301;
wire W4302;
wire W4303;
wire W4304;
wire W4305;
wire W4306;
wire W4307;
wire W4308;
wire W4309;
wire W4310;
wire W4311;
wire W4312;
wire W4313;
wire W4314;
wire W4315;
wire W4316;
wire W4317;
wire W4318;
wire W4319;
wire W4320;
wire W4321;
wire W4322;
wire W4323;
wire W4324;
wire W4325;
wire W4326;
wire W4327;
wire W4328;
wire W4329;
wire W4330;
wire W4331;
wire W4332;
wire W4333;
wire W4334;
wire W4335;
wire W4336;
wire W4337;
wire W4338;
wire W4339;
wire W4340;
wire W4341;
wire W4342;
wire W4343;
wire W4344;
wire W4345;
wire W4346;
wire W4347;
wire W4348;
wire W4349;
wire W4350;
wire W4351;
wire W4352;
wire W4353;
wire W4354;
wire W4355;
wire W4356;
wire W4357;
wire W4358;
wire W4359;
wire W4360;
wire W4361;
wire W4362;
wire W4363;
wire W4364;
wire W4365;
wire W4366;
wire W4367;
wire W4368;
wire W4369;
wire W4370;
wire W4371;
wire W4372;
wire W4373;
wire W4374;
wire W4375;
wire W4376;
wire W4377;
wire W4378;
wire W4379;
wire W4380;
wire W4381;
wire W4382;
wire W4383;
wire W4384;
wire W4385;
wire W4386;
wire W4387;
wire W4388;
wire W4389;
wire W4390;
wire W4391;
wire W4392;
wire W4393;
wire W4394;
wire W4395;
wire W4396;
wire W4397;
wire W4398;
wire W4399;
wire W4400;
wire W4401;
wire W4402;
wire W4403;
wire W4404;
wire W4405;
wire W4406;
wire W4407;
wire W4408;
wire W4409;
wire W4410;
wire W4411;
wire W4412;
wire W4413;
wire W4414;
wire W4415;
wire W4416;
wire W4417;
wire W4418;
wire W4419;
wire W4420;
wire W4421;
wire W4422;
wire W4423;
wire W4424;
wire W4425;
wire W4426;
wire W4427;
wire W4428;
wire W4429;
wire W4430;
wire W4431;
wire W4432;
wire W4433;
wire W4434;
wire W4435;
wire W4436;
wire W4437;
wire W4438;
wire W4439;
wire W4440;
wire W4441;
wire W4442;
wire W4443;
wire W4444;
wire W4445;
wire W4446;
wire W4447;
wire W4448;
wire W4449;
wire W4450;
wire W4451;
wire W4452;
wire W4453;
wire W4454;
wire W4455;
wire W4456;
wire W4457;
wire W4458;
wire W4459;
wire W4460;
wire W4461;
wire W4462;
wire W4463;
wire W4464;
wire W4465;
wire W4466;
wire W4467;
wire W4468;
wire W4469;
wire W4470;
wire W4471;
wire W4472;
wire W4473;
wire W4474;
wire W4475;
wire W4476;
wire W4477;
wire W4478;
wire W4479;
wire W4480;
wire W4481;
wire W4482;
wire W4483;
wire W4484;
wire W4485;
wire W4486;
wire W4487;
wire W4488;
wire W4489;
wire W4490;
wire W4491;
wire W4492;
wire W4493;
wire W4494;
wire W4495;
wire W4496;
wire W4497;
wire W4498;
wire W4499;
wire W4500;
wire W4501;
wire W4502;
wire W4503;
wire W4504;
wire W4505;
wire W4506;
wire W4507;
wire W4508;
wire W4509;
wire W4510;
wire W4511;
wire W4512;
wire W4513;
wire W4514;
wire W4515;
wire W4516;
wire W4517;
wire W4518;
wire W4519;
wire W4520;
wire W4521;
wire W4522;
wire W4523;
wire W4524;
wire W4525;
wire W4526;
wire W4527;
wire W4528;
wire W4529;
wire W4530;
wire W4531;
wire W4532;
wire W4533;
wire W4534;
wire W4535;
wire W4536;
wire W4537;
wire W4538;
wire W4539;
wire W4540;
wire W4541;
wire W4542;
wire W4543;
wire W4544;
wire W4545;
wire W4546;
wire W4547;
wire W4548;
wire W4549;
wire W4550;
wire W4551;
wire W4552;
wire W4553;
wire W4554;
wire W4555;
wire W4556;
wire W4557;
wire W4558;
wire W4559;
wire W4560;
wire W4561;
wire W4562;
wire W4563;
wire W4564;
wire W4565;
wire W4566;
wire W4567;
wire W4568;
wire W4569;
wire W4570;
wire W4571;
wire W4572;
wire W4573;
wire W4574;
wire W4575;
wire W4576;
wire W4577;
wire W4578;
wire W4579;
wire W4580;
wire W4581;
wire W4582;
wire W4583;
wire W4584;
wire W4585;
wire W4586;
wire W4587;
wire W4588;
wire W4589;
wire W4590;
wire W4591;
wire W4592;
wire W4593;
wire W4594;
wire W4595;
wire W4596;
wire W4597;
wire W4598;
wire W4599;
wire W4600;
wire W4601;
wire W4602;
wire W4603;
wire W4604;
wire W4605;
wire W4606;
wire W4607;
wire W4608;
wire W4609;
wire W4610;
wire W4611;
wire W4612;
wire W4613;
wire W4614;
wire W4615;
wire W4616;
wire W4617;
wire W4618;
wire W4619;
wire W4620;
wire W4621;
wire W4622;
wire W4623;
wire W4624;
wire W4625;
wire W4626;
wire W4627;
wire W4628;
wire W4629;
wire W4630;
wire W4631;
wire W4632;
wire W4633;
wire W4634;
wire W4635;
wire W4636;
wire W4637;
wire W4638;
wire W4639;
wire W4640;
wire W4641;
wire W4642;
wire W4643;
wire W4644;
wire W4645;
wire W4646;
wire W4647;
wire W4648;
wire W4649;
wire W4650;
wire W4651;
wire W4652;
wire W4653;
wire W4654;
wire W4655;
wire W4656;
wire W4657;
wire W4658;
wire W4659;
wire W4660;
wire W4661;
wire W4662;
wire W4663;
wire W4664;
wire W4665;
wire W4666;
wire W4667;
wire W4668;
wire W4669;
wire W4670;
wire W4671;
wire W4672;
wire W4673;
wire W4674;
wire W4675;
wire W4676;
wire W4677;
wire W4678;
wire W4679;
wire W4680;
wire W4681;
wire W4682;
wire W4683;
wire W4684;
wire W4685;
wire W4686;
wire W4687;
wire W4688;
wire W4689;
wire W4690;
wire W4691;
wire W4692;
wire W4693;
wire W4694;
wire W4695;
wire W4696;
wire W4697;
wire W4698;
wire W4699;
wire W4700;
wire W4701;
wire W4702;
wire W4703;
wire W4704;
wire W4705;
wire W4706;
wire W4707;
wire W4708;
wire W4709;
wire W4710;
wire W4711;
wire W4712;
wire W4713;
wire W4714;
wire W4715;
wire W4716;
wire W4717;
wire W4718;
wire W4719;
wire W4720;
wire W4721;
wire W4722;
wire W4723;
wire W4724;
wire W4725;
wire W4726;
wire W4727;
wire W4728;
wire W4729;
wire W4730;
wire W4731;
wire W4732;
wire W4733;
wire W4734;
wire W4735;
wire W4736;
wire W4737;
wire W4738;
wire W4739;
wire W4740;
wire W4741;
wire W4742;
wire W4743;
wire W4744;
wire W4745;
wire W4746;
wire W4747;
wire W4748;
wire W4749;
wire W4750;
wire W4751;
wire W4752;
wire W4753;
wire W4754;
wire W4755;
wire W4756;
wire W4757;
wire W4758;
wire W4759;
wire W4760;
wire W4761;
wire W4762;
wire W4763;
wire W4764;
wire W4765;
wire W4766;
wire W4767;
wire W4768;
wire W4769;
wire W4770;
wire W4771;
wire W4772;
wire W4773;
wire W4774;
wire W4775;
wire W4776;
wire W4777;
wire W4778;
wire W4779;
wire W4780;
wire W4781;
wire W4782;
wire W4783;
wire W4784;
wire W4785;
wire W4786;
wire W4787;
wire W4788;
wire W4789;
wire W4790;
wire W4791;
wire W4792;
wire W4793;
wire W4794;
wire W4795;
wire W4796;
wire W4797;
wire W4798;
wire W4799;
wire W4800;
wire W4801;
wire W4802;
wire W4803;
wire W4804;
wire W4805;
wire W4806;
wire W4807;
wire W4808;
wire W4809;
wire W4810;
wire W4811;
wire W4812;
wire W4813;
wire W4814;
wire W4815;
wire W4816;
wire W4817;
wire W4818;
wire W4819;
wire W4820;
wire W4821;
wire W4822;
wire W4823;
wire W4824;
wire W4825;
wire W4826;
wire W4827;
wire W4828;
wire W4829;
wire W4830;
wire W4831;
wire W4832;
wire W4833;
wire W4834;
wire W4835;
wire W4836;
wire W4837;
wire W4838;
wire W4839;
wire W4840;
wire W4841;
wire W4842;
wire W4843;
wire W4844;
wire W4845;
wire W4846;
wire W4847;
wire W4848;
wire W4849;
wire W4850;
wire W4851;
wire W4852;
wire W4853;
wire W4854;
wire W4855;
wire W4856;
wire W4857;
wire W4858;
wire W4859;
wire W4860;
wire W4861;
wire W4862;
wire W4863;
wire W4864;
wire W4865;
wire W4866;
wire W4867;
wire W4868;
wire W4869;
wire W4870;
wire W4871;
wire W4872;
wire W4873;
wire W4874;
wire W4875;
wire W4876;
wire W4877;
wire W4878;
wire W4879;
wire W4880;
wire W4881;
wire W4882;
wire W4883;
wire W4884;
wire W4885;
wire W4886;
wire W4887;
wire W4888;
wire W4889;
wire W4890;
wire W4891;
wire W4892;
wire W4893;
wire W4894;
wire W4895;
wire W4896;
wire W4897;
wire W4898;
wire W4899;
wire W4900;
wire W4901;
wire W4902;
wire W4903;
wire W4904;
wire W4905;
wire W4906;
wire W4907;
wire W4908;
wire W4909;
wire W4910;
wire W4911;
wire W4912;
wire W4913;
wire W4914;
wire W4915;
wire W4916;
wire W4917;
wire W4918;
wire W4919;
wire W4920;
wire W4921;
wire W4922;
wire W4923;
wire W4924;
wire W4925;
wire W4926;
wire W4927;
wire W4928;
wire W4929;
wire W4930;
wire W4931;
wire W4932;
wire W4933;
wire W4934;
wire W4935;
wire W4936;
wire W4937;
wire W4938;
wire W4939;
wire W4940;
wire W4941;
wire W4942;
wire W4943;
wire W4944;
wire W4945;
wire W4946;
wire W4947;
wire W4948;
wire W4949;
wire W4950;
wire W4951;
wire W4952;
wire W4953;
wire W4954;
wire W4955;
wire W4956;
wire W4957;
wire W4958;
wire W4959;
wire W4960;
wire W4961;
wire W4962;
wire W4963;
wire W4964;
wire W4965;
wire W4966;
wire W4967;
wire W4968;
wire W4969;
wire W4970;
wire W4971;
wire W4972;
wire W4973;
wire W4974;
wire W4975;
wire W4976;
wire W4977;
wire W4978;
wire W4979;
wire W4980;
wire W4981;
wire W4982;
wire W4983;
wire W4984;
wire W4985;
wire W4986;
wire W4987;
wire W4988;
wire W4989;
wire W4990;
wire W4991;
wire W4992;
wire W4993;
wire W4994;
wire W4995;
wire W4996;
wire W4997;
wire W4998;
wire W4999;
wire W5000;
wire W5001;
wire W5002;
wire W5003;
wire W5004;
wire W5005;
wire W5006;
wire W5007;
wire W5008;
wire W5009;
wire W5010;
wire W5011;
wire W5012;
wire W5013;
wire W5014;
wire W5015;
wire W5016;
wire W5017;
wire W5018;
wire W5019;
wire W5020;
wire W5021;
wire W5022;
wire W5023;
wire W5024;
wire W5025;
wire W5026;
wire W5027;
wire W5028;
wire W5029;
wire W5030;
wire W5031;
wire W5032;
wire W5033;
wire W5034;
wire W5035;
wire W5036;
wire W5037;
wire W5038;
wire W5039;
wire W5040;
wire W5041;
wire W5042;
wire W5043;
wire W5044;
wire W5045;
wire W5046;
wire W5047;
wire W5048;
wire W5049;
wire W5050;
wire W5051;
wire W5052;
wire W5053;
wire W5054;
wire W5055;
wire W5056;
wire W5057;
wire W5058;
wire W5059;
wire W5060;
wire W5061;
wire W5062;
wire W5063;
wire W5064;
wire W5065;
wire W5066;
wire W5067;
wire W5068;
wire W5069;
wire W5070;
wire W5071;
wire W5072;
wire W5073;
wire W5074;
wire W5075;
wire W5076;
wire W5077;
wire W5078;
wire W5079;
wire W5080;
wire W5081;
wire W5082;
wire W5083;
wire W5084;
wire W5085;
wire W5086;
wire W5087;
wire W5088;
wire W5089;
wire W5090;
wire W5091;
wire W5092;
wire W5093;
wire W5094;
wire W5095;
wire W5096;
wire W5097;
wire W5098;
wire W5099;
wire W5100;
wire W5101;
wire W5102;
wire W5103;
wire W5104;
wire W5105;
wire W5106;
wire W5107;
wire W5108;
wire W5109;
wire W5110;
wire W5111;
wire W5112;
wire W5113;
wire W5114;
wire W5115;
wire W5116;
wire W5117;
wire W5118;
wire W5119;
wire W5120;
wire W5121;
wire W5122;
wire W5123;
wire W5124;
wire W5125;
wire W5126;
wire W5127;
wire W5128;
wire W5129;
wire W5130;
wire W5131;
wire W5132;
wire W5133;
wire W5134;
wire W5135;
wire W5136;
wire W5137;
wire W5138;
wire W5139;
wire W5140;
wire W5141;
wire W5142;
wire W5143;
wire W5144;
wire W5145;
wire W5146;
wire W5147;
wire W5148;
wire W5149;
wire W5150;
wire W5151;
wire W5152;
wire W5153;
wire W5154;
wire W5155;
wire W5156;
wire W5157;
wire W5158;
wire W5159;
wire W5160;
wire W5161;
wire W5162;
wire W5163;
wire W5164;
wire W5165;
wire W5166;
wire W5167;
wire W5168;
wire W5169;
wire W5170;
wire W5171;
wire W5172;
wire W5173;
wire W5174;
wire W5175;
wire W5176;
wire W5177;
wire W5178;
wire W5179;
wire W5180;
wire W5181;
wire W5182;
wire W5183;
wire W5184;
wire W5185;
wire W5186;
wire W5187;
wire W5188;
wire W5189;
wire W5190;
wire W5191;
wire W5192;
wire W5193;
wire W5194;
wire W5195;
wire W5196;
wire W5197;
wire W5198;
wire W5199;
wire W5200;
wire W5201;
wire W5202;
wire W5203;
wire W5204;
wire W5205;
wire W5206;
wire W5207;
wire W5208;
wire W5209;
wire W5210;
wire W5211;
wire W5212;
wire W5213;
wire W5214;
wire W5215;
wire W5216;
wire W5217;
wire W5218;
wire W5219;
wire W5220;
wire W5221;
wire W5222;
wire W5223;
wire W5224;
wire W5225;
wire W5226;
wire W5227;
wire W5228;
wire W5229;
wire W5230;
wire W5231;
wire W5232;
wire W5233;
wire W5234;
wire W5235;
wire W5236;
wire W5237;
wire W5238;
wire W5239;
wire W5240;
wire W5241;
wire W5242;
wire W5243;
wire W5244;
wire W5245;
wire W5246;
wire W5247;
wire W5248;
wire W5249;
wire W5250;
wire W5251;
wire W5252;
wire W5253;
wire W5254;
wire W5255;
wire W5256;
wire W5257;
wire W5258;
wire W5259;
wire W5260;
wire W5261;
wire W5262;
wire W5263;
wire W5264;
wire W5265;
wire W5266;
wire W5267;
wire W5268;
wire W5269;
wire W5270;
wire W5271;
wire W5272;
wire W5273;
wire W5274;
wire W5275;
wire W5276;
wire W5277;
wire W5278;
wire W5279;
wire W5280;
wire W5281;
wire W5282;
wire W5283;
wire W5284;
wire W5285;
wire W5286;
wire W5287;
wire W5288;
wire W5289;
wire W5290;
wire W5291;
wire W5292;
wire W5293;
wire W5294;
wire W5295;
wire W5296;
wire W5297;
wire W5298;
wire W5299;
wire W5300;
wire W5301;
wire W5302;
wire W5303;
wire W5304;
wire W5305;
wire W5306;
wire W5307;
wire W5308;
wire W5309;
wire W5310;
wire W5311;
wire W5312;
wire W5313;
wire W5314;
wire W5315;
wire W5316;
wire W5317;
wire W5318;
wire W5319;
wire W5320;
wire W5321;
wire W5322;
wire W5323;
wire W5324;
wire W5325;
wire W5326;
wire W5327;
wire W5328;
wire W5329;
wire W5330;
wire W5331;
wire W5332;
wire W5333;
wire W5334;
wire W5335;
wire W5336;
wire W5337;
wire W5338;
wire W5339;
wire W5340;
wire W5341;
wire W5342;
wire W5343;
wire W5344;
wire W5345;
wire W5346;
wire W5347;
wire W5348;
wire W5349;
wire W5350;
wire W5351;
wire W5352;
wire W5353;
wire W5354;
wire W5355;
wire W5356;
wire W5357;
wire W5358;
wire W5359;
wire W5360;
wire W5361;
wire W5362;
wire W5363;
wire W5364;
wire W5365;
wire W5366;
wire W5367;
wire W5368;
wire W5369;
wire W5370;
wire W5371;
wire W5372;
wire W5373;
wire W5374;
wire W5375;
wire W5376;
wire W5377;
wire W5378;
wire W5379;
wire W5380;
wire W5381;
wire W5382;
wire W5383;
wire W5384;
wire W5385;
wire W5386;
wire W5387;
wire W5388;
wire W5389;
wire W5390;
wire W5391;
wire W5392;
wire W5393;
wire W5394;
wire W5395;
wire W5396;
wire W5397;
wire W5398;
wire W5399;
wire W5400;
wire W5401;
wire W5402;
wire W5403;
wire W5404;
wire W5405;
wire W5406;
wire W5407;
wire W5408;
wire W5409;
wire W5410;
wire W5411;
wire W5412;
wire W5413;
wire W5414;
wire W5415;
wire W5416;
wire W5417;
wire W5418;
wire W5419;
wire W5420;
wire W5421;
wire W5422;
wire W5423;
wire W5424;
wire W5425;
wire W5426;
wire W5427;
wire W5428;
wire W5429;
wire W5430;
wire W5431;
wire W5432;
wire W5433;
wire W5434;
wire W5435;
wire W5436;
wire W5437;
wire W5438;
wire W5439;
wire W5440;
wire W5441;
wire W5442;
wire W5443;
wire W5444;
wire W5445;
wire W5446;
wire W5447;
wire W5448;
wire W5449;
wire W5450;
wire W5451;
wire W5452;
wire W5453;
wire W5454;
wire W5455;
wire W5456;
wire W5457;
wire W5458;
wire W5459;
wire W5460;
wire W5461;
wire W5462;
wire W5463;
wire W5464;
wire W5465;
wire W5466;
wire W5467;
wire W5468;
wire W5469;
wire W5470;
wire W5471;
wire W5472;
wire W5473;
wire W5474;
wire W5475;
wire W5476;
wire W5477;
wire W5478;
wire W5479;
wire W5480;
wire W5481;
wire W5482;
wire W5483;
wire W5484;
wire W5485;
wire W5486;
wire W5487;
wire W5488;
wire W5489;
wire W5490;
wire W5491;
wire W5492;
wire W5493;
wire W5494;
wire W5495;
wire W5496;
wire W5497;
wire W5498;
wire W5499;
wire W5500;
wire W5501;
wire W5502;
wire W5503;
wire W5504;
wire W5505;
wire W5506;
wire W5507;
wire W5508;
wire W5509;
wire W5510;
wire W5511;
wire W5512;
wire W5513;
wire W5514;
wire W5515;
wire W5516;
wire W5517;
wire W5518;
wire W5519;
wire W5520;
wire W5521;
wire W5522;
wire W5523;
wire W5524;
wire W5525;
wire W5526;
wire W5527;
wire W5528;
wire W5529;
wire W5530;
wire W5531;
wire W5532;
wire W5533;
wire W5534;
wire W5535;
wire W5536;
wire W5537;
wire W5538;
wire W5539;
wire W5540;
wire W5541;
wire W5542;
wire W5543;
wire W5544;
wire W5545;
wire W5546;
wire W5547;
wire W5548;
wire W5549;
wire W5550;
wire W5551;
wire W5552;
wire W5553;
wire W5554;
wire W5555;
wire W5556;
wire W5557;
wire W5558;
wire W5559;
wire W5560;
wire W5561;
wire W5562;
wire W5563;
wire W5564;
wire W5565;
wire W5566;
wire W5567;
wire W5568;
wire W5569;
wire W5570;
wire W5571;
wire W5572;
wire W5573;
wire W5574;
wire W5575;
wire W5576;
wire W5577;
wire W5578;
wire W5579;
wire W5580;
wire W5581;
wire W5582;
wire W5583;
wire W5584;
wire W5585;
wire W5586;
wire W5587;
wire W5588;
wire W5589;
wire W5590;
wire W5591;
wire W5592;
wire W5593;
wire W5594;
wire W5595;
wire W5596;
wire W5597;
wire W5598;
wire W5599;
wire W5600;
wire W5601;
wire W5602;
wire W5603;
wire W5604;
wire W5605;
wire W5606;
wire W5607;
wire W5608;
wire W5609;
wire W5610;
wire W5611;
wire W5612;
wire W5613;
wire W5614;
wire W5615;
wire W5616;
wire W5617;
wire W5618;
wire W5619;
wire W5620;
wire W5621;
wire W5622;
wire W5623;
wire W5624;
wire W5625;
wire W5626;
wire W5627;
wire W5628;
wire W5629;
wire W5630;
wire W5631;
wire W5632;
wire W5633;
wire W5634;
wire W5635;
wire W5636;
wire W5637;
wire W5638;
wire W5639;
wire W5640;
wire W5641;
wire W5642;
wire W5643;
wire W5644;
wire W5645;
wire W5646;
wire W5647;
wire W5648;
wire W5649;
wire W5650;
wire W5651;
wire W5652;
wire W5653;
wire W5654;
wire W5655;
wire W5656;
wire W5657;
wire W5658;
wire W5659;
wire W5660;
wire W5661;
wire W5662;
wire W5663;
wire W5664;
wire W5665;
wire W5666;
wire W5667;
wire W5668;
wire W5669;
wire W5670;
wire W5671;
wire W5672;
wire W5673;
wire W5674;
wire W5675;
wire W5676;
wire W5677;
wire W5678;
wire W5679;
wire W5680;
wire W5681;
wire W5682;
wire W5683;
wire W5684;
wire W5685;
wire W5686;
wire W5687;
wire W5688;
wire W5689;
wire W5690;
wire W5691;
wire W5692;
wire W5693;
wire W5694;
wire W5695;
wire W5696;
wire W5697;
wire W5698;
wire W5699;
wire W5700;
wire W5701;
wire W5702;
wire W5703;
wire W5704;
wire W5705;
wire W5706;
wire W5707;
wire W5708;
wire W5709;
wire W5710;
wire W5711;
wire W5712;
wire W5713;
wire W5714;
wire W5715;
wire W5716;
wire W5717;
wire W5718;
wire W5719;
wire W5720;
wire W5721;
wire W5722;
wire W5723;
wire W5724;
wire W5725;
wire W5726;
wire W5727;
wire W5728;
wire W5729;
wire W5730;
wire W5731;
wire W5732;
wire W5733;
wire W5734;
wire W5735;
wire W5736;
wire W5737;
wire W5738;
wire W5739;
wire W5740;
wire W5741;
wire W5742;
wire W5743;
wire W5744;
wire W5745;
wire W5746;
wire W5747;
wire W5748;
wire W5749;
wire W5750;
wire W5751;
wire W5752;
wire W5753;
wire W5754;
wire W5755;
wire W5756;
wire W5757;
wire W5758;
wire W5759;
wire W5760;
wire W5761;
wire W5762;
wire W5763;
wire W5764;
wire W5765;
wire W5766;
wire W5767;
wire W5768;
wire W5769;
wire W5770;
wire W5771;
wire W5772;
wire W5773;
wire W5774;
wire W5775;
wire W5776;
wire W5777;
wire W5778;
wire W5779;
wire W5780;
wire W5781;
wire W5782;
wire W5783;
wire W5784;
wire W5785;
wire W5786;
wire W5787;
wire W5788;
wire W5789;
wire W5790;
wire W5791;
wire W5792;
wire W5793;
wire W5794;
wire W5795;
wire W5796;
wire W5797;
wire W5798;
wire W5799;
wire W5800;
wire W5801;
wire W5802;
wire W5803;
wire W5804;
wire W5805;
wire W5806;
wire W5807;
wire W5808;
wire W5809;
wire W5810;
wire W5811;
wire W5812;
wire W5813;
wire W5814;
wire W5815;
wire W5816;
wire W5817;
wire W5818;
wire W5819;
wire W5820;
wire W5821;
wire W5822;
wire W5823;
wire W5824;
wire W5825;
wire W5826;
wire W5827;
wire W5828;
wire W5829;
wire W5830;
wire W5831;
wire W5832;
wire W5833;
wire W5834;
wire W5835;
wire W5836;
wire W5837;
wire W5838;
wire W5839;
wire W5840;
wire W5841;
wire W5842;
wire W5843;
wire W5844;
wire W5845;
wire W5846;
wire W5847;
wire W5848;
wire W5849;
wire W5850;
wire W5851;
wire W5852;
wire W5853;
wire W5854;
wire W5855;
wire W5856;
wire W5857;
wire W5858;
wire W5859;
wire W5860;
wire W5861;
wire W5862;
wire W5863;
wire W5864;
wire W5865;
wire W5866;
wire W5867;
wire W5868;
wire W5869;
wire W5870;
wire W5871;
wire W5872;
wire W5873;
wire W5874;
wire W5875;
wire W5876;
wire W5877;
wire W5878;
wire W5879;
wire W5880;
wire W5881;
wire W5882;
wire W5883;
wire W5884;
wire W5885;
wire W5886;
wire W5887;
wire W5888;
wire W5889;
wire W5890;
wire W5891;
wire W5892;
wire W5893;
wire W5894;
wire W5895;
wire W5896;
wire W5897;
wire W5898;
wire W5899;
wire W5900;
wire W5901;
wire W5902;
wire W5903;
wire W5904;
wire W5905;
wire W5906;
wire W5907;
wire W5908;
wire W5909;
wire W5910;
wire W5911;
wire W5912;
wire W5913;
wire W5914;
wire W5915;
wire W5916;
wire W5917;
wire W5918;
wire W5919;
wire W5920;
wire W5921;
wire W5922;
wire W5923;
wire W5924;
wire W5925;
wire W5926;
wire W5927;
wire W5928;
wire W5929;
wire W5930;
wire W5931;
wire W5932;
wire W5933;
wire W5934;
wire W5935;
wire W5936;
wire W5937;
wire W5938;
wire W5939;
wire W5940;
wire W5941;
wire W5942;
wire W5943;
wire W5944;
wire W5945;
wire W5946;
wire W5947;
wire W5948;
wire W5949;
wire W5950;
wire W5951;
wire W5952;
wire W5953;
wire W5954;
wire W5955;
wire W5956;
wire W5957;
wire W5958;
wire W5959;
wire W5960;
wire W5961;
wire W5962;
wire W5963;
wire W5964;
wire W5965;
wire W5966;
wire W5967;
wire W5968;
wire W5969;
wire W5970;
wire W5971;
wire W5972;
wire W5973;
wire W5974;
wire W5975;
wire W5976;
wire W5977;
wire W5978;
wire W5979;
wire W5980;
wire W5981;
wire W5982;
wire W5983;
wire W5984;
wire W5985;
wire W5986;
wire W5987;
wire W5988;
wire W5989;
wire W5990;
wire W5991;
wire W5992;
wire W5993;
wire W5994;
wire W5995;
wire W5996;
wire W5997;
wire W5998;
wire W5999;
wire W6000;
wire W6001;
wire W6002;
wire W6003;
wire W6004;
wire W6005;
wire W6006;
wire W6007;
wire W6008;
wire W6009;
wire W6010;
wire W6011;
wire W6012;
wire W6013;
wire W6014;
wire W6015;
wire W6016;
wire W6017;
wire W6018;
wire W6019;
wire W6020;
wire W6021;
wire W6022;
wire W6023;
wire W6024;
wire W6025;
wire W6026;
wire W6027;
wire W6028;
wire W6029;
wire W6030;
wire W6031;
wire W6032;
wire W6033;
wire W6034;
wire W6035;
wire W6036;
wire W6037;
wire W6038;
wire W6039;
wire W6040;
wire W6041;
wire W6042;
wire W6043;
wire W6044;
wire W6045;
wire W6046;
wire W6047;
wire W6048;
wire W6049;
wire W6050;
wire W6051;
wire W6052;
wire W6053;
wire W6054;
wire W6055;
wire W6056;
wire W6057;
wire W6058;
wire W6059;
wire W6060;
wire W6061;
wire W6062;
wire W6063;
wire W6064;
wire W6065;
wire W6066;
wire W6067;
wire W6068;
wire W6069;
wire W6070;
wire W6071;
wire W6072;
wire W6073;
wire W6074;
wire W6075;
wire W6076;
wire W6077;
wire W6078;
wire W6079;
wire W6080;
wire W6081;
wire W6082;
wire W6083;
wire W6084;
wire W6085;
wire W6086;
wire W6087;
wire W6088;
wire W6089;
wire W6090;
wire W6091;
wire W6092;
wire W6093;
wire W6094;
wire W6095;
wire W6096;
wire W6097;
wire W6098;
wire W6099;
wire W6100;
wire W6101;
wire W6102;
wire W6103;
wire W6104;
wire W6105;
wire W6106;
wire W6107;
wire W6108;
wire W6109;
wire W6110;
wire W6111;
wire W6112;
wire W6113;
wire W6114;
wire W6115;
wire W6116;
wire W6117;
wire W6118;
wire W6119;
wire W6120;
wire W6121;
wire W6122;
wire W6123;
wire W6124;
wire W6125;
wire W6126;
wire W6127;
wire W6128;
wire W6129;
wire W6130;
wire W6131;
wire W6132;
wire W6133;
wire W6134;
wire W6135;
wire W6136;
wire W6137;
wire W6138;
wire W6139;
wire W6140;
wire W6141;
wire W6142;
wire W6143;
wire W6144;
wire W6145;
wire W6146;
wire W6147;
wire W6148;
wire W6149;
wire W6150;
wire W6151;
wire W6152;
wire W6153;
wire W6154;
wire W6155;
wire W6156;
wire W6157;
wire W6158;
wire W6159;
wire W6160;
wire W6161;
wire W6162;
wire W6163;
wire W6164;
wire W6165;
wire W6166;
wire W6167;
wire W6168;
wire W6169;
wire W6170;
wire W6171;
wire W6172;
wire W6173;
wire W6174;
wire W6175;
wire W6176;
wire W6177;
wire W6178;
wire W6179;
wire W6180;
wire W6181;
wire W6182;
wire W6183;
wire W6184;
wire W6185;
wire W6186;
wire W6187;
wire W6188;
wire W6189;
wire W6190;
wire W6191;
wire W6192;
wire W6193;
wire W6194;
wire W6195;
wire W6196;
wire W6197;
wire W6198;
wire W6199;
wire W6200;
wire W6201;
wire W6202;
wire W6203;
wire W6204;
wire W6205;
wire W6206;
wire W6207;
wire W6208;
wire W6209;
wire W6210;
wire W6211;
wire W6212;
wire W6213;
wire W6214;
wire W6215;
wire W6216;
wire W6217;
wire W6218;
wire W6219;
wire W6220;
wire W6221;
wire W6222;
wire W6223;
wire W6224;
wire W6225;
wire W6226;
wire W6227;
wire W6228;
wire W6229;
wire W6230;
wire W6231;
wire W6232;
wire W6233;
wire W6234;
wire W6235;
wire W6236;
wire W6237;
wire W6238;
wire W6239;
wire W6240;
wire W6241;
wire W6242;
wire W6243;
wire W6244;
wire W6245;
wire W6246;
wire W6247;
wire W6248;
wire W6249;
wire W6250;
wire W6251;
wire W6252;
wire W6253;
wire W6254;
wire W6255;
wire W6256;
wire W6257;
wire W6258;
wire W6259;
wire W6260;
wire W6261;
wire W6262;
wire W6263;
wire W6264;
wire W6265;
wire W6266;
wire W6267;
wire W6268;
wire W6269;
wire W6270;
wire W6271;
wire W6272;
wire W6273;
wire W6274;
wire W6275;
wire W6276;
wire W6277;
wire W6278;
wire W6279;
wire W6280;
wire W6281;
wire W6282;
wire W6283;
wire W6284;
wire W6285;
wire W6286;
wire W6287;
wire W6288;
wire W6289;
wire W6290;
wire W6291;
wire W6292;
wire W6293;
wire W6294;
wire W6295;
wire W6296;
wire W6297;
wire W6298;
wire W6299;
wire W6300;
wire W6301;
wire W6302;
wire W6303;
wire W6304;
wire W6305;
wire W6306;
wire W6307;
wire W6308;
wire W6309;
wire W6310;
wire W6311;
wire W6312;
wire W6313;
wire W6314;
wire W6315;
wire W6316;
wire W6317;
wire W6318;
wire W6319;
wire W6320;
wire W6321;
wire W6322;
wire W6323;
wire W6324;
wire W6325;
wire W6326;
wire W6327;
wire W6328;
wire W6329;
wire W6330;
wire W6331;
wire W6332;
wire W6333;
wire W6334;
wire W6335;
wire W6336;
wire W6337;
wire W6338;
wire W6339;
wire W6340;
wire W6341;
wire W6342;
wire W6343;
wire W6344;
wire W6345;
wire W6346;
wire W6347;
wire W6348;
wire W6349;
wire W6350;
wire W6351;
wire W6352;
wire W6353;
wire W6354;
wire W6355;
wire W6356;
wire W6357;
wire W6358;
wire W6359;
wire W6360;
wire W6361;
wire W6362;
wire W6363;
wire W6364;
wire W6365;
wire W6366;
wire W6367;
wire W6368;
wire W6369;
wire W6370;
wire W6371;
wire W6372;
wire W6373;
wire W6374;
wire W6375;
wire W6376;
wire W6377;
wire W6378;
wire W6379;
wire W6380;
wire W6381;
wire W6382;
wire W6383;
wire W6384;
wire W6385;
wire W6386;
wire W6387;
wire W6388;
wire W6389;
wire W6390;
wire W6391;
wire W6392;
wire W6393;
wire W6394;
wire W6395;
wire W6396;
wire W6397;
wire W6398;
wire W6399;
wire W6400;
wire W6401;
wire W6402;
wire W6403;
wire W6404;
wire W6405;
wire W6406;
wire W6407;
wire W6408;
wire W6409;
wire W6410;
wire W6411;
wire W6412;
wire W6413;
wire W6414;
wire W6415;
wire W6416;
wire W6417;
wire W6418;
wire W6419;
wire W6420;
wire W6421;
wire W6422;
wire W6423;
wire W6424;
wire W6425;
wire W6426;
wire W6427;
wire W6428;
wire W6429;
wire W6430;
wire W6431;
wire W6432;
wire W6433;
wire W6434;
wire W6435;
wire W6436;
wire W6437;
wire W6438;
wire W6439;
wire W6440;
wire W6441;
wire W6442;
wire W6443;
wire W6444;
wire W6445;
wire W6446;
wire W6447;
wire W6448;
wire W6449;
wire W6450;
wire W6451;
wire W6452;
wire W6453;
wire W6454;
wire W6455;
wire W6456;
wire W6457;
wire W6458;
wire W6459;
wire W6460;
wire W6461;
wire W6462;
wire W6463;
wire W6464;
wire W6465;
wire W6466;
wire W6467;
wire W6468;
wire W6469;
wire W6470;
wire W6471;
wire W6472;
wire W6473;
wire W6474;
wire W6475;
wire W6476;
wire W6477;
wire W6478;
wire W6479;
wire W6480;
wire W6481;
wire W6482;
wire W6483;
wire W6484;
wire W6485;
wire W6486;
wire W6487;
wire W6488;
wire W6489;
wire W6490;
wire W6491;
wire W6492;
wire W6493;
wire W6494;
wire W6495;
wire W6496;
wire W6497;
wire W6498;
wire W6499;
wire W6500;
wire W6501;
wire W6502;
wire W6503;
wire W6504;
wire W6505;
wire W6506;
wire W6507;
wire W6508;
wire W6509;
wire W6510;
wire W6511;
wire W6512;
wire W6513;
wire W6514;
wire W6515;
wire W6516;
wire W6517;
wire W6518;
wire W6519;
wire W6520;
wire W6521;
wire W6522;
wire W6523;
wire W6524;
wire W6525;
wire W6526;
wire W6527;
wire W6528;
wire W6529;
wire W6530;
wire W6531;
wire W6532;
wire W6533;
wire W6534;
wire W6535;
wire W6536;
wire W6537;
wire W6538;
wire W6539;
wire W6540;
wire W6541;
wire W6542;
wire W6543;
wire W6544;
wire W6545;
wire W6546;
wire W6547;
wire W6548;
wire W6549;
wire W6550;
wire W6551;
wire W6552;
wire W6553;
wire W6554;
wire W6555;
wire W6556;
wire W6557;
wire W6558;
wire W6559;
wire W6560;
wire W6561;
wire W6562;
wire W6563;
wire W6564;
wire W6565;
wire W6566;
wire W6567;
wire W6568;
wire W6569;
wire W6570;
wire W6571;
wire W6572;
wire W6573;
wire W6574;
wire W6575;
wire W6576;
wire W6577;
wire W6578;
wire W6579;
wire W6580;
wire W6581;
wire W6582;
wire W6583;
wire W6584;
wire W6585;
wire W6586;
wire W6587;
wire W6588;
wire W6589;
wire W6590;
wire W6591;
wire W6592;
wire W6593;
wire W6594;
wire W6595;
wire W6596;
wire W6597;
wire W6598;
wire W6599;
wire W6600;
wire W6601;
wire W6602;
wire W6603;
wire W6604;
wire W6605;
wire W6606;
wire W6607;
wire W6608;
wire W6609;
wire W6610;
wire W6611;
wire W6612;
wire W6613;
wire W6614;
wire W6615;
wire W6616;
wire W6617;
wire W6618;
wire W6619;
wire W6620;
wire W6621;
wire W6622;
wire W6623;
wire W6624;
wire W6625;
wire W6626;
wire W6627;
wire W6628;
wire W6629;
wire W6630;
wire W6631;
wire W6632;
wire W6633;
wire W6634;
wire W6635;
wire W6636;
wire W6637;
wire W6638;
wire W6639;
wire W6640;
wire W6641;
wire W6642;
wire W6643;
wire W6644;
wire W6645;
wire W6646;
wire W6647;
wire W6648;
wire W6649;
wire W6650;
wire W6651;
wire W6652;
wire W6653;
wire W6654;
wire W6655;
wire W6656;
wire W6657;
wire W6658;
wire W6659;
wire W6660;
wire W6661;
wire W6662;
wire W6663;
wire W6664;
wire W6665;
wire W6666;
wire W6667;
wire W6668;
wire W6669;
wire W6670;
wire W6671;
wire W6672;
wire W6673;
wire W6674;
wire W6675;
wire W6676;
wire W6677;
wire W6678;
wire W6679;
wire W6680;
wire W6681;
wire W6682;
wire W6683;
wire W6684;
wire W6685;
wire W6686;
wire W6687;
wire W6688;
wire W6689;
wire W6690;
wire W6691;
wire W6692;
wire W6693;
wire W6694;
wire W6695;
wire W6696;
wire W6697;
wire W6698;
wire W6699;
wire W6700;
wire W6701;
wire W6702;
wire W6703;
wire W6704;
wire W6705;
wire W6706;
wire W6707;
wire W6708;
wire W6709;
wire W6710;
wire W6711;
wire W6712;
wire W6713;
wire W6714;
wire W6715;
wire W6716;
wire W6717;
wire W6718;
wire W6719;
wire W6720;
wire W6721;
wire W6722;
wire W6723;
wire W6724;
wire W6725;
wire W6726;
wire W6727;
wire W6728;
wire W6729;
wire W6730;
wire W6731;
wire W6732;
wire W6733;
wire W6734;
wire W6735;
wire W6736;
wire W6737;
wire W6738;
wire W6739;
wire W6740;
wire W6741;
wire W6742;
wire W6743;
wire W6744;
wire W6745;
wire W6746;
wire W6747;
wire W6748;
wire W6749;
wire W6750;
wire W6751;
wire W6752;
wire W6753;
wire W6754;
wire W6755;
wire W6756;
wire W6757;
wire W6758;
wire W6759;
wire W6760;
wire W6761;
wire W6762;
wire W6763;
wire W6764;
wire W6765;
wire W6766;
wire W6767;
wire W6768;
wire W6769;
wire W6770;
wire W6771;
wire W6772;
wire W6773;
wire W6774;
wire W6775;
wire W6776;
wire W6777;
wire W6778;
wire W6779;
wire W6780;
wire W6781;
wire W6782;
wire W6783;
wire W6784;
wire W6785;
wire W6786;
wire W6787;
wire W6788;
wire W6789;
wire W6790;
wire W6791;
wire W6792;
wire W6793;
wire W6794;
wire W6795;
wire W6796;
wire W6797;
wire W6798;
wire W6799;
wire W6800;
wire W6801;
wire W6802;
wire W6803;
wire W6804;
wire W6805;
wire W6806;
wire W6807;
wire W6808;
wire W6809;
wire W6810;
wire W6811;
wire W6812;
wire W6813;
wire W6814;
wire W6815;
wire W6816;
wire W6817;
wire W6818;
wire W6819;
wire W6820;
wire W6821;
wire W6822;
wire W6823;
wire W6824;
wire W6825;
wire W6826;
wire W6827;
wire W6828;
wire W6829;
wire W6830;
wire W6831;
wire W6832;
wire W6833;
wire W6834;
wire W6835;
wire W6836;
wire W6837;
wire W6838;
wire W6839;
wire W6840;
wire W6841;
wire W6842;
wire W6843;
wire W6844;
wire W6845;
wire W6846;
wire W6847;
wire W6848;
wire W6849;
wire W6850;
wire W6851;
wire W6852;
wire W6853;
wire W6854;
wire W6855;
wire W6856;
wire W6857;
wire W6858;
wire W6859;
wire W6860;
wire W6861;
wire W6862;
wire W6863;
wire W6864;
wire W6865;
wire W6866;
wire W6867;
wire W6868;
wire W6869;
wire W6870;
wire W6871;
wire W6872;
wire W6873;
wire W6874;
wire W6875;
wire W6876;
wire W6877;
wire W6878;
wire W6879;
wire W6880;
wire W6881;
wire W6882;
wire W6883;
wire W6884;
wire W6885;
wire W6886;
wire W6887;
wire W6888;
wire W6889;
wire W6890;
wire W6891;
wire W6892;
wire W6893;
wire W6894;
wire W6895;
wire W6896;
wire W6897;
wire W6898;
wire W6899;
wire W6900;
wire W6901;
wire W6902;
wire W6903;
wire W6904;
wire W6905;
wire W6906;
wire W6907;
wire W6908;
wire W6909;
wire W6910;
wire W6911;
wire W6912;
wire W6913;
wire W6914;
wire W6915;
wire W6916;
wire W6917;
wire W6918;
wire W6919;
wire W6920;
wire W6921;
wire W6922;
wire W6923;
wire W6924;
wire W6925;
wire W6926;
wire W6927;
wire W6928;
wire W6929;
wire W6930;
wire W6931;
wire W6932;
wire W6933;
wire W6934;
wire W6935;
wire W6936;
wire W6937;
wire W6938;
wire W6939;
wire W6940;
wire W6941;
wire W6942;
wire W6943;
wire W6944;
wire W6945;
wire W6946;
wire W6947;
wire W6948;
wire W6949;
wire W6950;
wire W6951;
wire W6952;
wire W6953;
wire W6954;
wire W6955;
wire W6956;
wire W6957;
wire W6958;
wire W6959;
wire W6960;
wire W6961;
wire W6962;
wire W6963;
wire W6964;
wire W6965;
wire W6966;
wire W6967;
wire W6968;
wire W6969;
wire W6970;
wire W6971;
wire W6972;
wire W6973;
wire W6974;
wire W6975;
wire W6976;
wire W6977;
wire W6978;
wire W6979;
wire W6980;
wire W6981;
wire W6982;
wire W6983;
wire W6984;
wire W6985;
wire W6986;
wire W6987;
wire W6988;
wire W6989;
wire W6990;
wire W6991;
wire W6992;
wire W6993;
wire W6994;
wire W6995;
wire W6996;
wire W6997;
wire W6998;
wire W6999;
wire W7000;
wire W7001;
wire W7002;
wire W7003;
wire W7004;
wire W7005;
wire W7006;
wire W7007;
wire W7008;
wire W7009;
wire W7010;
wire W7011;
wire W7012;
wire W7013;
wire W7014;
wire W7015;
wire W7016;
wire W7017;
wire W7018;
wire W7019;
wire W7020;
wire W7021;
wire W7022;
wire W7023;
wire W7024;
wire W7025;
wire W7026;
wire W7027;
wire W7028;
wire W7029;
wire W7030;
wire W7031;
wire W7032;
wire W7033;
wire W7034;
wire W7035;
wire W7036;
wire W7037;
wire W7038;
wire W7039;
wire W7040;
wire W7041;
wire W7042;
wire W7043;
wire W7044;
wire W7045;
wire W7046;
wire W7047;
wire W7048;
wire W7049;
wire W7050;
wire W7051;
wire W7052;
wire W7053;
wire W7054;
wire W7055;
wire W7056;
wire W7057;
wire W7058;
wire W7059;
wire W7060;
wire W7061;
wire W7062;
wire W7063;
wire W7064;
wire W7065;
wire W7066;
wire W7067;
wire W7068;
wire W7069;
wire W7070;
wire W7071;
wire W7072;
wire W7073;
wire W7074;
wire W7075;
wire W7076;
wire W7077;
wire W7078;
wire W7079;
wire W7080;
wire W7081;
wire W7082;
wire W7083;
wire W7084;
wire W7085;
wire W7086;
wire W7087;
wire W7088;
wire W7089;
wire W7090;
wire W7091;
wire W7092;
wire W7093;
wire W7094;
wire W7095;
wire W7096;
wire W7097;
wire W7098;
wire W7099;
wire W7100;
wire W7101;
wire W7102;
wire W7103;
wire W7104;
wire W7105;
wire W7106;
wire W7107;
wire W7108;
wire W7109;
wire W7110;
wire W7111;
wire W7112;
wire W7113;
wire W7114;
wire W7115;
wire W7116;
wire W7117;
wire W7118;
wire W7119;
wire W7120;
wire W7121;
wire W7122;
wire W7123;
wire W7124;
wire W7125;
wire W7126;
wire W7127;
wire W7128;
wire W7129;
wire W7130;
wire W7131;
wire W7132;
wire W7133;
wire W7134;
wire W7135;
wire W7136;
wire W7137;
wire W7138;
wire W7139;
wire W7140;
wire W7141;
wire W7142;
wire W7143;
wire W7144;
wire W7145;
wire W7146;
wire W7147;
wire W7148;
wire W7149;
wire W7150;
wire W7151;
wire W7152;
wire W7153;
wire W7154;
wire W7155;
wire W7156;
wire W7157;
wire W7158;
wire W7159;
wire W7160;
wire W7161;
wire W7162;
wire W7163;
wire W7164;
wire W7165;
wire W7166;
wire W7167;
wire W7168;
wire W7169;
wire W7170;
wire W7171;
wire W7172;
wire W7173;
wire W7174;
wire W7175;
wire W7176;
wire W7177;
wire W7178;
wire W7179;
wire W7180;
wire W7181;
wire W7182;
wire W7183;
wire W7184;
wire W7185;
wire W7186;
wire W7187;
wire W7188;
wire W7189;
wire W7190;
wire W7191;
wire W7192;
wire W7193;
wire W7194;
wire W7195;
wire W7196;
wire W7197;
wire W7198;
wire W7199;
wire W7200;
wire W7201;
wire W7202;
wire W7203;
wire W7204;
wire W7205;
wire W7206;
wire W7207;
wire W7208;
wire W7209;
wire W7210;
wire W7211;
wire W7212;
wire W7213;
wire W7214;
wire W7215;
wire W7216;
wire W7217;
wire W7218;
wire W7219;
wire W7220;
wire W7221;
wire W7222;
wire W7223;
wire W7224;
wire W7225;
wire W7226;
wire W7227;
wire W7228;
wire W7229;
wire W7230;
wire W7231;
wire W7232;
wire W7233;
wire W7234;
wire W7235;
wire W7236;
wire W7237;
wire W7238;
wire W7239;
wire W7240;
wire W7241;
wire W7242;
wire W7243;
wire W7244;
wire W7245;
wire W7246;
wire W7247;
wire W7248;
wire W7249;
wire W7250;
wire W7251;
wire W7252;
wire W7253;
wire W7254;
wire W7255;
wire W7256;
wire W7257;
wire W7258;
wire W7259;
wire W7260;
wire W7261;
wire W7262;
wire W7263;
wire W7264;
wire W7265;
wire W7266;
wire W7267;
wire W7268;
wire W7269;
wire W7270;
wire W7271;
wire W7272;
wire W7273;
wire W7274;
wire W7275;
wire W7276;
wire W7277;
wire W7278;
wire W7279;
wire W7280;
wire W7281;
wire W7282;
wire W7283;
wire W7284;
wire W7285;
wire W7286;
wire W7287;
wire W7288;
wire W7289;
wire W7290;
wire W7291;
wire W7292;
wire W7293;
wire W7294;
wire W7295;
wire W7296;
wire W7297;
wire W7298;
wire W7299;
wire W7300;
wire W7301;
wire W7302;
wire W7303;
wire W7304;
wire W7305;
wire W7306;
wire W7307;
wire W7308;
wire W7309;
wire W7310;
wire W7311;
wire W7312;
wire W7313;
wire W7314;
wire W7315;
wire W7316;
wire W7317;
wire W7318;
wire W7319;
wire W7320;
wire W7321;
wire W7322;
wire W7323;
wire W7324;
wire W7325;
wire W7326;
wire W7327;
wire W7328;
wire W7329;
wire W7330;
wire W7331;
wire W7332;
wire W7333;
wire W7334;
wire W7335;
wire W7336;
wire W7337;
wire W7338;
wire W7339;
wire W7340;
wire W7341;
wire W7342;
wire W7343;
wire W7344;
wire W7345;
wire W7346;
wire W7347;
wire W7348;
wire W7349;
wire W7350;
wire W7351;
wire W7352;
wire W7353;
wire W7354;
wire W7355;
wire W7356;
wire W7357;
wire W7358;
wire W7359;
wire W7360;
wire W7361;
wire W7362;
wire W7363;
wire W7364;
wire W7365;
wire W7366;
wire W7367;
wire W7368;
wire W7369;
wire W7370;
wire W7371;
wire W7372;
wire W7373;
wire W7374;
wire W7375;
wire W7376;
wire W7377;
wire W7378;
wire W7379;
wire W7380;
wire W7381;
wire W7382;
wire W7383;
wire W7384;
wire W7385;
wire W7386;
wire W7387;
wire W7388;
wire W7389;
wire W7390;
wire W7391;
wire W7392;
wire W7393;
wire W7394;
wire W7395;
wire W7396;
wire W7397;
wire W7398;
wire W7399;
wire W7400;
wire W7401;
wire W7402;
wire W7403;
wire W7404;
wire W7405;
wire W7406;
wire W7407;
wire W7408;
wire W7409;
wire W7410;
wire W7411;
wire W7412;
wire W7413;
wire W7414;
wire W7415;
wire W7416;
wire W7417;
wire W7418;
wire W7419;
wire W7420;
wire W7421;
wire W7422;
wire W7423;
wire W7424;
wire W7425;
wire W7426;
wire W7427;
wire W7428;
wire W7429;
wire W7430;
wire W7431;
wire W7432;
wire W7433;
wire W7434;
wire W7435;
wire W7436;
wire W7437;
wire W7438;
wire W7439;
wire W7440;
wire W7441;
wire W7442;
wire W7443;
wire W7444;
wire W7445;
wire W7446;
wire W7447;
wire W7448;
wire W7449;
wire W7450;
wire W7451;
wire W7452;
wire W7453;
wire W7454;
wire W7455;
wire W7456;
wire W7457;
wire W7458;
wire W7459;
wire W7460;
wire W7461;
wire W7462;
wire W7463;
wire W7464;
wire W7465;
wire W7466;
wire W7467;
wire W7468;
wire W7469;
wire W7470;
wire W7471;
wire W7472;
wire W7473;
wire W7474;
wire W7475;
wire W7476;
wire W7477;
wire W7478;
wire W7479;
wire W7480;
wire W7481;
wire W7482;
wire W7483;
wire W7484;
wire W7485;
wire W7486;
wire W7487;
wire W7488;
wire W7489;
wire W7490;
wire W7491;
wire W7492;
wire W7493;
wire W7494;
wire W7495;
wire W7496;
wire W7497;
wire W7498;
wire W7499;
wire W7500;
wire W7501;
wire W7502;
wire W7503;
wire W7504;
wire W7505;
wire W7506;
wire W7507;
wire W7508;
wire W7509;
wire W7510;
wire W7511;
wire W7512;
wire W7513;
wire W7514;
wire W7515;
wire W7516;
wire W7517;
wire W7518;
wire W7519;
wire W7520;
wire W7521;
wire W7522;
wire W7523;
wire W7524;
wire W7525;
wire W7526;
wire W7527;
wire W7528;
wire W7529;
wire W7530;
wire W7531;
wire W7532;
wire W7533;
wire W7534;
wire W7535;
wire W7536;
wire W7537;
wire W7538;
wire W7539;
wire W7540;
wire W7541;
wire W7542;
wire W7543;
wire W7544;
wire W7545;
wire W7546;
wire W7547;
wire W7548;
wire W7549;
wire W7550;
wire W7551;
wire W7552;
wire W7553;
wire W7554;
wire W7555;
wire W7556;
wire W7557;
wire W7558;
wire W7559;
wire W7560;
wire W7561;
wire W7562;
wire W7563;
wire W7564;
wire W7565;
wire W7566;
wire W7567;
wire W7568;
wire W7569;
wire W7570;
wire W7571;
wire W7572;
wire W7573;
wire W7574;
wire W7575;
wire W7576;
wire W7577;
wire W7578;
wire W7579;
wire W7580;
wire W7581;
wire W7582;
wire W7583;
wire W7584;
wire W7585;
wire W7586;
wire W7587;
wire W7588;
wire W7589;
wire W7590;
wire W7591;
wire W7592;
wire W7593;
wire W7594;
wire W7595;
wire W7596;
wire W7597;
wire W7598;
wire W7599;
wire W7600;
wire W7601;
wire W7602;
wire W7603;
wire W7604;
wire W7605;
wire W7606;
wire W7607;
wire W7608;
wire W7609;
wire W7610;
wire W7611;
wire W7612;
wire W7613;
wire W7614;
wire W7615;
wire W7616;
wire W7617;
wire W7618;
wire W7619;
wire W7620;
wire W7621;
wire W7622;
wire W7623;
wire W7624;
wire W7625;
wire W7626;
wire W7627;
wire W7628;
wire W7629;
wire W7630;
wire W7631;
wire W7632;
wire W7633;
wire W7634;
wire W7635;
wire W7636;
wire W7637;
wire W7638;
wire W7639;
wire W7640;
wire W7641;
wire W7642;
wire W7643;
wire W7644;
wire W7645;
wire W7646;
wire W7647;
wire W7648;
wire W7649;
wire W7650;
wire W7651;
wire W7652;
wire W7653;
wire W7654;
wire W7655;
wire W7656;
wire W7657;
wire W7658;
wire W7659;
wire W7660;
wire W7661;
wire W7662;
wire W7663;
wire W7664;
wire W7665;
wire W7666;
wire W7667;
wire W7668;
wire W7669;
wire W7670;
wire W7671;
wire W7672;
wire W7673;
wire W7674;
wire W7675;
wire W7676;
wire W7677;
wire W7678;
wire W7679;
wire W7680;
wire W7681;
wire W7682;
wire W7683;
wire W7684;
wire W7685;
wire W7686;
wire W7687;
wire W7688;
wire W7689;
wire W7690;
wire W7691;
wire W7692;
wire W7693;
wire W7694;
wire W7695;
wire W7696;
wire W7697;
wire W7698;
wire W7699;
wire W7700;
wire W7701;
wire W7702;
wire W7703;
wire W7704;
wire W7705;
wire W7706;
wire W7707;
wire W7708;
wire W7709;
wire W7710;
wire W7711;
wire W7712;
wire W7713;
wire W7714;
wire W7715;
wire W7716;
wire W7717;
wire W7718;
wire W7719;
wire W7720;
wire W7721;
wire W7722;
wire W7723;
wire W7724;
wire W7725;
wire W7726;
wire W7727;
wire W7728;
wire W7729;
wire W7730;
wire W7731;
wire W7732;
wire W7733;
wire W7734;
wire W7735;
wire W7736;
wire W7737;
wire W7738;
wire W7739;
wire W7740;
wire W7741;
wire W7742;
wire W7743;
wire W7744;
wire W7745;
wire W7746;
wire W7747;
wire W7748;
wire W7749;
wire W7750;
wire W7751;
wire W7752;
wire W7753;
wire W7754;
wire W7755;
wire W7756;
wire W7757;
wire W7758;
wire W7759;
wire W7760;
wire W7761;
wire W7762;
wire W7763;
wire W7764;
wire W7765;
wire W7766;
wire W7767;
wire W7768;
wire W7769;
wire W7770;
wire W7771;
wire W7772;
wire W7773;
wire W7774;
wire W7775;
wire W7776;
wire W7777;
wire W7778;
wire W7779;
wire W7780;
wire W7781;
wire W7782;
wire W7783;
wire W7784;
wire W7785;
wire W7786;
wire W7787;
wire W7788;
wire W7789;
wire W7790;
wire W7791;
wire W7792;
wire W7793;
wire W7794;
wire W7795;
wire W7796;
wire W7797;
wire W7798;
wire W7799;
wire W7800;
wire W7801;
wire W7802;
wire W7803;
wire W7804;
wire W7805;
wire W7806;
wire W7807;
wire W7808;
wire W7809;
wire W7810;
wire W7811;
wire W7812;
wire W7813;
wire W7814;
wire W7815;
wire W7816;
wire W7817;
wire W7818;
wire W7819;
wire W7820;
wire W7821;
wire W7822;
wire W7823;
wire W7824;
wire W7825;
wire W7826;
wire W7827;
wire W7828;
wire W7829;
wire W7830;
wire W7831;
wire W7832;
wire W7833;
wire W7834;
wire W7835;
wire W7836;
wire W7837;
wire W7838;
wire W7839;
wire W7840;
wire W7841;
wire W7842;
wire W7843;
wire W7844;
wire W7845;
wire W7846;
wire W7847;
wire W7848;
wire W7849;
wire W7850;
wire W7851;
wire W7852;
wire W7853;
wire W7854;
wire W7855;
wire W7856;
wire W7857;
wire W7858;
wire W7859;
wire W7860;
wire W7861;
wire W7862;
wire W7863;
wire W7864;
wire W7865;
wire W7866;
wire W7867;
wire W7868;
wire W7869;
wire W7870;
wire W7871;
wire W7872;
wire W7873;
wire W7874;
wire W7875;
wire W7876;
wire W7877;
wire W7878;
wire W7879;
wire W7880;
wire W7881;
wire W7882;
wire W7883;
wire W7884;
wire W7885;
wire W7886;
wire W7887;
wire W7888;
wire W7889;
wire W7890;
wire W7891;
wire W7892;
wire W7893;
wire W7894;
wire W7895;
wire W7896;
wire W7897;
wire W7898;
wire W7899;
wire W7900;
wire W7901;
wire W7902;
wire W7903;
wire W7904;
wire W7905;
wire W7906;
wire W7907;
wire W7908;
wire W7909;
wire W7910;
wire W7911;
wire W7912;
wire W7913;
wire W7914;
wire W7915;
wire W7916;
wire W7917;
wire W7918;
wire W7919;
wire W7920;
wire W7921;
wire W7922;
wire W7923;
wire W7924;
wire W7925;
wire W7926;
wire W7927;
wire W7928;
wire W7929;
wire W7930;
wire W7931;
wire W7932;
wire W7933;
wire W7934;
wire W7935;
wire W7936;
wire W7937;
wire W7938;
wire W7939;
wire W7940;
wire W7941;
wire W7942;
wire W7943;
wire W7944;
wire W7945;
wire W7946;
wire W7947;
wire W7948;
wire W7949;
wire W7950;
wire W7951;
wire W7952;
wire W7953;
wire W7954;
wire W7955;
wire W7956;
wire W7957;
wire W7958;
wire W7959;
wire W7960;
wire W7961;
wire W7962;
wire W7963;
wire W7964;
wire W7965;
wire W7966;
wire W7967;
wire W7968;
wire W7969;
wire W7970;
wire W7971;
wire W7972;
wire W7973;
wire W7974;
wire W7975;
wire W7976;
wire W7977;
wire W7978;
wire W7979;
wire W7980;
wire W7981;
wire W7982;
wire W7983;
wire W7984;
wire W7985;
wire W7986;
wire W7987;
wire W7988;
wire W7989;
wire W7990;
wire W7991;
wire W7992;
wire W7993;
wire W7994;
wire W7995;
wire W7996;
wire W7997;
wire W7998;
wire W7999;
wire W8000;
wire W8001;
wire W8002;
wire W8003;
wire W8004;
wire W8005;
wire W8006;
wire W8007;
wire W8008;
wire W8009;
wire W8010;
wire W8011;
wire W8012;
wire W8013;
wire W8014;
wire W8015;
wire W8016;
wire W8017;
wire W8018;
wire W8019;
wire W8020;
wire W8021;
wire W8022;
wire W8023;
wire W8024;
wire W8025;
wire W8026;
wire W8027;
wire W8028;
wire W8029;
wire W8030;
wire W8031;
wire W8032;
wire W8033;
wire W8034;
wire W8035;
wire W8036;
wire W8037;
wire W8038;
wire W8039;
wire W8040;
wire W8041;
wire W8042;
wire W8043;
wire W8044;
wire W8045;
wire W8046;
wire W8047;
wire W8048;
wire W8049;
wire W8050;
wire W8051;
wire W8052;
wire W8053;
wire W8054;
wire W8055;
wire W8056;
wire W8057;
wire W8058;
wire W8059;
wire W8060;
wire W8061;
wire W8062;
wire W8063;
wire W8064;
wire W8065;
wire W8066;
wire W8067;
wire W8068;
wire W8069;
wire W8070;
wire W8071;
wire W8072;
wire W8073;
wire W8074;
wire W8075;
wire W8076;
wire W8077;
wire W8078;
wire W8079;
wire W8080;
wire W8081;
wire W8082;
wire W8083;
wire W8084;
wire W8085;
wire W8086;
wire W8087;
wire W8088;
wire W8089;
wire W8090;
wire W8091;
wire W8092;
wire W8093;
wire W8094;
wire W8095;
wire W8096;
wire W8097;
wire W8098;
wire W8099;
wire W8100;
wire W8101;
wire W8102;
wire W8103;
wire W8104;
wire W8105;
wire W8106;
wire W8107;
wire W8108;
wire W8109;
wire W8110;
wire W8111;
wire W8112;
wire W8113;
wire W8114;
wire W8115;
wire W8116;
wire W8117;
wire W8118;
wire W8119;
wire W8120;
wire W8121;
wire W8122;
wire W8123;
wire W8124;
wire W8125;
wire W8126;
wire W8127;
wire W8128;
wire W8129;
wire W8130;
wire W8131;
wire W8132;
wire W8133;
wire W8134;
wire W8135;
wire W8136;
wire W8137;
wire W8138;
wire W8139;
wire W8140;
wire W8141;
wire W8142;
wire W8143;
wire W8144;
wire W8145;
wire W8146;
wire W8147;
wire W8148;
wire W8149;
wire W8150;
wire W8151;
wire W8152;
wire W8153;
wire W8154;
wire W8155;
wire W8156;
wire W8157;
wire W8158;
wire W8159;
wire W8160;
wire W8161;
wire W8162;
wire W8163;
wire W8164;
wire W8165;
wire W8166;
wire W8167;
wire W8168;
wire W8169;
wire W8170;
wire W8171;
wire W8172;
wire W8173;
wire W8174;
wire W8175;
wire W8176;
wire W8177;
wire W8178;
wire W8179;
wire W8180;
wire W8181;
wire W8182;
wire W8183;
wire W8184;
wire W8185;
wire W8186;
wire W8187;
wire W8188;
wire W8189;
wire W8190;
wire W8191;
wire W8192;
wire W8193;
wire W8194;
wire W8195;
wire W8196;
wire W8197;
wire W8198;
wire W8199;
wire W8200;
wire W8201;
wire W8202;
wire W8203;
wire W8204;
wire W8205;
wire W8206;
wire W8207;
wire W8208;
wire W8209;
wire W8210;
wire W8211;
wire W8212;
wire W8213;
wire W8214;
wire W8215;
wire W8216;
wire W8217;
wire W8218;
wire W8219;
wire W8220;
wire W8221;
wire W8222;
wire W8223;
wire W8224;
wire W8225;
wire W8226;
wire W8227;
wire W8228;
wire W8229;
wire W8230;
wire W8231;
wire W8232;
wire W8233;
wire W8234;
wire W8235;
wire W8236;
wire W8237;
wire W8238;
wire W8239;
wire W8240;
wire W8241;
wire W8242;
wire W8243;
wire W8244;
wire W8245;
wire W8246;
wire W8247;
wire W8248;
wire W8249;
wire W8250;
wire W8251;
wire W8252;
wire W8253;
wire W8254;
wire W8255;
wire W8256;
wire W8257;
wire W8258;
wire W8259;
wire W8260;
wire W8261;
wire W8262;
wire W8263;
wire W8264;
wire W8265;
wire W8266;
wire W8267;
wire W8268;
wire W8269;
wire W8270;
wire W8271;
wire W8272;
wire W8273;
wire W8274;
wire W8275;
wire W8276;
wire W8277;
wire W8278;
wire W8279;
wire W8280;
wire W8281;
wire W8282;
wire W8283;
wire W8284;
wire W8285;
wire W8286;
wire W8287;
wire W8288;
wire W8289;
wire W8290;
wire W8291;
wire W8292;
wire W8293;
wire W8294;
wire W8295;
wire W8296;
wire W8297;
wire W8298;
wire W8299;
wire W8300;
wire W8301;
wire W8302;
wire W8303;
wire W8304;
wire W8305;
wire W8306;
wire W8307;
wire W8308;
wire W8309;
wire W8310;
wire W8311;
wire W8312;
wire W8313;
wire W8314;
wire W8315;
wire W8316;
wire W8317;
wire W8318;
wire W8319;
wire W8320;
wire W8321;
wire W8322;
wire W8323;
wire W8324;
wire W8325;
wire W8326;
wire W8327;
wire W8328;
wire W8329;
wire W8330;
wire W8331;
wire W8332;
wire W8333;
wire W8334;
wire W8335;
wire W8336;
wire W8337;
wire W8338;
wire W8339;
wire W8340;
wire W8341;
wire W8342;
wire W8343;
wire W8344;
wire W8345;
wire W8346;
wire W8347;
wire W8348;
wire W8349;
wire W8350;
wire W8351;
wire W8352;
wire W8353;
wire W8354;
wire W8355;
wire W8356;
wire W8357;
wire W8358;
wire W8359;
wire W8360;
wire W8361;
wire W8362;
wire W8363;
wire W8364;
wire W8365;
wire W8366;
wire W8367;
wire W8368;
wire W8369;
wire W8370;
wire W8371;
wire W8372;
wire W8373;
wire W8374;
wire W8375;
wire W8376;
wire W8377;
wire W8378;
wire W8379;
wire W8380;
wire W8381;
wire W8382;
wire W8383;
wire W8384;
wire W8385;
wire W8386;
wire W8387;
wire W8388;
wire W8389;
wire W8390;
wire W8391;
wire W8392;
wire W8393;
wire W8394;
wire W8395;
wire W8396;
wire W8397;
wire W8398;
wire W8399;
wire W8400;
wire W8401;
wire W8402;
wire W8403;
wire W8404;
wire W8405;
wire W8406;
wire W8407;
wire W8408;
wire W8409;
wire W8410;
wire W8411;
wire W8412;
wire W8413;
wire W8414;
wire W8415;
wire W8416;
wire W8417;
wire W8418;
wire W8419;
wire W8420;
wire W8421;
wire W8422;
wire W8423;
wire W8424;
wire W8425;
wire W8426;
wire W8427;
wire W8428;
wire W8429;
wire W8430;
wire W8431;
wire W8432;
wire W8433;
wire W8434;
wire W8435;
wire W8436;
wire W8437;
wire W8438;
wire W8439;
wire W8440;
wire W8441;
wire W8442;
wire W8443;
wire W8444;
wire W8445;
wire W8446;
wire W8447;
wire W8448;
wire W8449;
wire W8450;
wire W8451;
wire W8452;
wire W8453;
wire W8454;
wire W8455;
wire W8456;
wire W8457;
wire W8458;
wire W8459;
wire W8460;
wire W8461;
wire W8462;
wire W8463;
wire W8464;
wire W8465;
wire W8466;
wire W8467;
wire W8468;
wire W8469;
wire W8470;
wire W8471;
wire W8472;
wire W8473;
wire W8474;
wire W8475;
wire W8476;
wire W8477;
wire W8478;
wire W8479;
wire W8480;
wire W8481;
wire W8482;
wire W8483;
wire W8484;
wire W8485;
wire W8486;
wire W8487;
wire W8488;
wire W8489;
wire W8490;
wire W8491;
wire W8492;
wire W8493;
wire W8494;
wire W8495;
wire W8496;
wire W8497;
wire W8498;
wire W8499;
wire W8500;
wire W8501;
wire W8502;
wire W8503;
wire W8504;
wire W8505;
wire W8506;
wire W8507;
wire W8508;
wire W8509;
wire W8510;
wire W8511;
wire W8512;
wire W8513;
wire W8514;
wire W8515;
wire W8516;
wire W8517;
wire W8518;
wire W8519;
wire W8520;
wire W8521;
wire W8522;
wire W8523;
wire W8524;
wire W8525;
wire W8526;
wire W8527;
wire W8528;
wire W8529;
wire W8530;
wire W8531;
wire W8532;
wire W8533;
wire W8534;
wire W8535;
wire W8536;
wire W8537;
wire W8538;
wire W8539;
wire W8540;
wire W8541;
wire W8542;
wire W8543;
wire W8544;
wire W8545;
wire W8546;
wire W8547;
wire W8548;
wire W8549;
wire W8550;
wire W8551;
wire W8552;
wire W8553;
wire W8554;
wire W8555;
wire W8556;
wire W8557;
wire W8558;
wire W8559;
wire W8560;
wire W8561;
wire W8562;
wire W8563;
wire W8564;
wire W8565;
wire W8566;
wire W8567;
wire W8568;
wire W8569;
wire W8570;
wire W8571;
wire W8572;
wire W8573;
wire W8574;
wire W8575;
wire W8576;
wire W8577;
wire W8578;
wire W8579;
wire W8580;
wire W8581;
wire W8582;
wire W8583;
wire W8584;
wire W8585;
wire W8586;
wire W8587;
wire W8588;
wire W8589;
wire W8590;
wire W8591;
wire W8592;
wire W8593;
wire W8594;
wire W8595;
wire W8596;
wire W8597;
wire W8598;
wire W8599;
wire W8600;
wire W8601;
wire W8602;
wire W8603;
wire W8604;
wire W8605;
wire W8606;
wire W8607;
wire W8608;
wire W8609;
wire W8610;
wire W8611;
wire W8612;
wire W8613;
wire W8614;
wire W8615;
wire W8616;
wire W8617;
wire W8618;
wire W8619;
wire W8620;
wire W8621;
wire W8622;
wire W8623;
wire W8624;
wire W8625;
wire W8626;
wire W8627;
wire W8628;
wire W8629;
wire W8630;
wire W8631;
wire W8632;
wire W8633;
wire W8634;
wire W8635;
wire W8636;
wire W8637;
wire W8638;
wire W8639;
wire W8640;
wire W8641;
wire W8642;
wire W8643;
wire W8644;
wire W8645;
wire W8646;
wire W8647;
wire W8648;
wire W8649;
wire W8650;
wire W8651;
wire W8652;
wire W8653;
wire W8654;
wire W8655;
wire W8656;
wire W8657;
wire W8658;
wire W8659;
wire W8660;
wire W8661;
wire W8662;
wire W8663;
wire W8664;
wire W8665;
wire W8666;
wire W8667;
wire W8668;
wire W8669;
wire W8670;
wire W8671;
wire W8672;
wire W8673;
wire W8674;
wire W8675;
wire W8676;
wire W8677;
wire W8678;
wire W8679;
wire W8680;
wire W8681;
wire W8682;
wire W8683;
wire W8684;
wire W8685;
wire W8686;
wire W8687;
wire W8688;
wire W8689;
wire W8690;
wire W8691;
wire W8692;
wire W8693;
wire W8694;
wire W8695;
wire W8696;
wire W8697;
wire W8698;
wire W8699;
wire W8700;
wire W8701;
wire W8702;
wire W8703;
wire W8704;
wire W8705;
wire W8706;
wire W8707;
wire W8708;
wire W8709;
wire W8710;
wire W8711;
wire W8712;
wire W8713;
wire W8714;
wire W8715;
wire W8716;
wire W8717;
wire W8718;
wire W8719;
wire W8720;
wire W8721;
wire W8722;
wire W8723;
wire W8724;
wire W8725;
wire W8726;
wire W8727;
wire W8728;
wire W8729;
wire W8730;
wire W8731;
wire W8732;
wire W8733;
wire W8734;
wire W8735;
wire W8736;
wire W8737;
wire W8738;
wire W8739;
wire W8740;
wire W8741;
wire W8742;
wire W8743;
wire W8744;
wire W8745;
wire W8746;
wire W8747;
wire W8748;
wire W8749;
wire W8750;
wire W8751;
wire W8752;
wire W8753;
wire W8754;
wire W8755;
wire W8756;
wire W8757;
wire W8758;
wire W8759;
wire W8760;
wire W8761;
wire W8762;
wire W8763;
wire W8764;
wire W8765;
wire W8766;
wire W8767;
wire W8768;
wire W8769;
wire W8770;
wire W8771;
wire W8772;
wire W8773;
wire W8774;
wire W8775;
wire W8776;
wire W8777;
wire W8778;
wire W8779;
wire W8780;
wire W8781;
wire W8782;
wire W8783;
wire W8784;
wire W8785;
wire W8786;
wire W8787;
wire W8788;
wire W8789;
wire W8790;
wire W8791;
wire W8792;
wire W8793;
wire W8794;
wire W8795;
wire W8796;
wire W8797;
wire W8798;
wire W8799;
wire W8800;
wire W8801;
wire W8802;
wire W8803;
wire W8804;
wire W8805;
wire W8806;
wire W8807;
wire W8808;
wire W8809;
wire W8810;
wire W8811;
wire W8812;
wire W8813;
wire W8814;
wire W8815;
wire W8816;
wire W8817;
wire W8818;
wire W8819;
wire W8820;
wire W8821;
wire W8822;
wire W8823;
wire W8824;
wire W8825;
wire W8826;
wire W8827;
wire W8828;
wire W8829;
wire W8830;
wire W8831;
wire W8832;
wire W8833;
wire W8834;
wire W8835;
wire W8836;
wire W8837;
wire W8838;
wire W8839;
wire W8840;
wire W8841;
wire W8842;
wire W8843;
wire W8844;
wire W8845;
wire W8846;
wire W8847;
wire W8848;
wire W8849;
wire W8850;
wire W8851;
wire W8852;
wire W8853;
wire W8854;
wire W8855;
wire W8856;
wire W8857;
wire W8858;
wire W8859;
wire W8860;
wire W8861;
wire W8862;
wire W8863;
wire W8864;
wire W8865;
wire W8866;
wire W8867;
wire W8868;
wire W8869;
wire W8870;
wire W8871;
wire W8872;
wire W8873;
wire W8874;
wire W8875;
wire W8876;
wire W8877;
wire W8878;
wire W8879;
wire W8880;
wire W8881;
wire W8882;
wire W8883;
wire W8884;
wire W8885;
wire W8886;
wire W8887;
wire W8888;
wire W8889;
wire W8890;
wire W8891;
wire W8892;
wire W8893;
wire W8894;
wire W8895;
wire W8896;
wire W8897;
wire W8898;
wire W8899;
wire W8900;
wire W8901;
wire W8902;
wire W8903;
wire W8904;
wire W8905;
wire W8906;
wire W8907;
wire W8908;
wire W8909;
wire W8910;
wire W8911;
wire W8912;
wire W8913;
wire W8914;
wire W8915;
wire W8916;
wire W8917;
wire W8918;
wire W8919;
wire W8920;
wire W8921;
wire W8922;
wire W8923;
wire W8924;
wire W8925;
wire W8926;
wire W8927;
wire W8928;
wire W8929;
wire W8930;
wire W8931;
wire W8932;
wire W8933;
wire W8934;
wire W8935;
wire W8936;
wire W8937;
wire W8938;
wire W8939;
wire W8940;
wire W8941;
wire W8942;
wire W8943;
wire W8944;
wire W8945;
wire W8946;
wire W8947;
wire W8948;
wire W8949;
wire W8950;
wire W8951;
wire W8952;
wire W8953;
wire W8954;
wire W8955;
wire W8956;
wire W8957;
wire W8958;
wire W8959;
wire W8960;
wire W8961;
wire W8962;
wire W8963;
wire W8964;
wire W8965;
wire W8966;
wire W8967;
wire W8968;
wire W8969;
wire W8970;
wire W8971;
wire W8972;
wire W8973;
wire W8974;
wire W8975;
wire W8976;
wire W8977;
wire W8978;
wire W8979;
wire W8980;
wire W8981;
wire W8982;
wire W8983;
wire W8984;
wire W8985;
wire W8986;
wire W8987;
wire W8988;
wire W8989;
wire W8990;
wire W8991;
wire W8992;
wire W8993;
wire W8994;
wire W8995;
wire W8996;
wire W8997;
wire W8998;
wire W8999;
wire W9000;
wire W9001;
wire W9002;
wire W9003;
wire W9004;
wire W9005;
wire W9006;
wire W9007;
wire W9008;
wire W9009;
wire W9010;
wire W9011;
wire W9012;
wire W9013;
wire W9014;
wire W9015;
wire W9016;
wire W9017;
wire W9018;
wire W9019;
wire W9020;
wire W9021;
wire W9022;
wire W9023;
wire W9024;
wire W9025;
wire W9026;
wire W9027;
wire W9028;
wire W9029;
wire W9030;
wire W9031;
wire W9032;
wire W9033;
wire W9034;
wire W9035;
wire W9036;
wire W9037;
wire W9038;
wire W9039;
wire W9040;
wire W9041;
wire W9042;
wire W9043;
wire W9044;
wire W9045;
wire W9046;
wire W9047;
wire W9048;
wire W9049;
wire W9050;
wire W9051;
wire W9052;
wire W9053;
wire W9054;
wire W9055;
wire W9056;
wire W9057;
wire W9058;
wire W9059;
wire W9060;
wire W9061;
wire W9062;
wire W9063;
wire W9064;
wire W9065;
wire W9066;
wire W9067;
wire W9068;
wire W9069;
wire W9070;
wire W9071;
wire W9072;
wire W9073;
wire W9074;
wire W9075;
wire W9076;
wire W9077;
wire W9078;
wire W9079;
wire W9080;
wire W9081;
wire W9082;
wire W9083;
wire W9084;
wire W9085;
wire W9086;
wire W9087;
wire W9088;
wire W9089;
wire W9090;
wire W9091;
wire W9092;
wire W9093;
wire W9094;
wire W9095;
wire W9096;
wire W9097;
wire W9098;
wire W9099;
wire W9100;
wire W9101;
wire W9102;
wire W9103;
wire W9104;
wire W9105;
wire W9106;
wire W9107;
wire W9108;
wire W9109;
wire W9110;
wire W9111;
wire W9112;
wire W9113;
wire W9114;
wire W9115;
wire W9116;
wire W9117;
wire W9118;
wire W9119;
wire W9120;
wire W9121;
wire W9122;
wire W9123;
wire W9124;
wire W9125;
wire W9126;
wire W9127;
wire W9128;
wire W9129;
wire W9130;
wire W9131;
wire W9132;
wire W9133;
wire W9134;
wire W9135;
wire W9136;
wire W9137;
wire W9138;
wire W9139;
wire W9140;
wire W9141;
wire W9142;
wire W9143;
wire W9144;
wire W9145;
wire W9146;
wire W9147;
wire W9148;
wire W9149;
wire W9150;
wire W9151;
wire W9152;
wire W9153;
wire W9154;
wire W9155;
wire W9156;
wire W9157;
wire W9158;
wire W9159;
wire W9160;
wire W9161;
wire W9162;
wire W9163;
wire W9164;
wire W9165;
wire W9166;
wire W9167;
wire W9168;
wire W9169;
wire W9170;
wire W9171;
wire W9172;
wire W9173;
wire W9174;
wire W9175;
wire W9176;
wire W9177;
wire W9178;
wire W9179;
wire W9180;
wire W9181;
wire W9182;
wire W9183;
wire W9184;
wire W9185;
wire W9186;
wire W9187;
wire W9188;
wire W9189;
wire W9190;
wire W9191;
wire W9192;
wire W9193;
wire W9194;
wire W9195;
wire W9196;
wire W9197;
wire W9198;
wire W9199;
wire W9200;
wire W9201;
wire W9202;
wire W9203;
wire W9204;
wire W9205;
wire W9206;
wire W9207;
wire W9208;
wire W9209;
wire W9210;
wire W9211;
wire W9212;
wire W9213;
wire W9214;
wire W9215;
wire W9216;
wire W9217;
wire W9218;
wire W9219;
wire W9220;
wire W9221;
wire W9222;
wire W9223;
wire W9224;
wire W9225;
wire W9226;
wire W9227;
wire W9228;
wire W9229;
wire W9230;
wire W9231;
wire W9232;
wire W9233;
wire W9234;
wire W9235;
wire W9236;
wire W9237;
wire W9238;
wire W9239;
wire W9240;
wire W9241;
wire W9242;
wire W9243;
wire W9244;
wire W9245;
wire W9246;
wire W9247;
wire W9248;
wire W9249;
wire W9250;
wire W9251;
wire W9252;
wire W9253;
wire W9254;
wire W9255;
wire W9256;
wire W9257;
wire W9258;
wire W9259;
wire W9260;
wire W9261;
wire W9262;
wire W9263;
wire W9264;
wire W9265;
wire W9266;
wire W9267;
wire W9268;
wire W9269;
wire W9270;
wire W9271;
wire W9272;
wire W9273;
wire W9274;
wire W9275;
wire W9276;
wire W9277;
wire W9278;
wire W9279;
wire W9280;
wire W9281;
wire W9282;
wire W9283;
wire W9284;
wire W9285;
wire W9286;
wire W9287;
wire W9288;
wire W9289;
wire W9290;
wire W9291;
wire W9292;
wire W9293;
wire W9294;
wire W9295;
wire W9296;
wire W9297;
wire W9298;
wire W9299;
wire W9300;
wire W9301;
wire W9302;
wire W9303;
wire W9304;
wire W9305;
wire W9306;
wire W9307;
wire W9308;
wire W9309;
wire W9310;
wire W9311;
wire W9312;
wire W9313;
wire W9314;
wire W9315;
wire W9316;
wire W9317;
wire W9318;
wire W9319;
wire W9320;
wire W9321;
wire W9322;
wire W9323;
wire W9324;
wire W9325;
wire W9326;
wire W9327;
wire W9328;
wire W9329;
wire W9330;
wire W9331;
wire W9332;
wire W9333;
wire W9334;
wire W9335;
wire W9336;
wire W9337;
wire W9338;
wire W9339;
wire W9340;
wire W9341;
wire W9342;
wire W9343;
wire W9344;
wire W9345;
wire W9346;
wire W9347;
wire W9348;
wire W9349;
wire W9350;
wire W9351;
wire W9352;
wire W9353;
wire W9354;
wire W9355;
wire W9356;
wire W9357;
wire W9358;
wire W9359;
wire W9360;
wire W9361;
wire W9362;
wire W9363;
wire W9364;
wire W9365;
wire W9366;
wire W9367;
wire W9368;
wire W9369;
wire W9370;
wire W9371;
wire W9372;
wire W9373;
wire W9374;
wire W9375;
wire W9376;
wire W9377;
wire W9378;
wire W9379;
wire W9380;
wire W9381;
wire W9382;
wire W9383;
wire W9384;
wire W9385;
wire W9386;
wire W9387;
wire W9388;
wire W9389;
wire W9390;
wire W9391;
wire W9392;
wire W9393;
wire W9394;
wire W9395;
wire W9396;
wire W9397;
wire W9398;
wire W9399;
wire W9400;
wire W9401;
wire W9402;
wire W9403;
wire W9404;
wire W9405;
wire W9406;
wire W9407;
wire W9408;
wire W9409;
wire W9410;
wire W9411;
wire W9412;
wire W9413;
wire W9414;
wire W9415;
wire W9416;
wire W9417;
wire W9418;
wire W9419;
wire W9420;
wire W9421;
wire W9422;
wire W9423;
wire W9424;
wire W9425;
wire W9426;
wire W9427;
wire W9428;
wire W9429;
wire W9430;
wire W9431;
wire W9432;
wire W9433;
wire W9434;
wire W9435;
wire W9436;
wire W9437;
wire W9438;
wire W9439;
wire W9440;
wire W9441;
wire W9442;
wire W9443;
wire W9444;
wire W9445;
wire W9446;
wire W9447;
wire W9448;
wire W9449;
wire W9450;
wire W9451;
wire W9452;
wire W9453;
wire W9454;
wire W9455;
wire W9456;
wire W9457;
wire W9458;
wire W9459;
wire W9460;
wire W9461;
wire W9462;
wire W9463;
wire W9464;
wire W9465;
wire W9466;
wire W9467;
wire W9468;
wire W9469;
wire W9470;
wire W9471;
wire W9472;
wire W9473;
wire W9474;
wire W9475;
wire W9476;
wire W9477;
wire W9478;
wire W9479;
wire W9480;
wire W9481;
wire W9482;
wire W9483;
wire W9484;
wire W9485;
wire W9486;
wire W9487;
wire W9488;
wire W9489;
wire W9490;
wire W9491;
wire W9492;
wire W9493;
wire W9494;
wire W9495;
wire W9496;
wire W9497;
wire W9498;
wire W9499;
wire W9500;
wire W9501;
wire W9502;
wire W9503;
wire W9504;
wire W9505;
wire W9506;
wire W9507;
wire W9508;
wire W9509;
wire W9510;
wire W9511;
wire W9512;
wire W9513;
wire W9514;
wire W9515;
wire W9516;
wire W9517;
wire W9518;
wire W9519;
wire W9520;
wire W9521;
wire W9522;
wire W9523;
wire W9524;
wire W9525;
wire W9526;
wire W9527;
wire W9528;
wire W9529;
wire W9530;
wire W9531;
wire W9532;
wire W9533;
wire W9534;
wire W9535;
wire W9536;
wire W9537;
wire W9538;
wire W9539;
wire W9540;
wire W9541;
wire W9542;
wire W9543;
wire W9544;
wire W9545;
wire W9546;
wire W9547;
wire W9548;
wire W9549;
wire W9550;
wire W9551;
wire W9552;
wire W9553;
wire W9554;
wire W9555;
wire W9556;
wire W9557;
wire W9558;
wire W9559;
wire W9560;
wire W9561;
wire W9562;
wire W9563;
wire W9564;
wire W9565;
wire W9566;
wire W9567;
wire W9568;
wire W9569;
wire W9570;
wire W9571;
wire W9572;
wire W9573;
wire W9574;
wire W9575;
wire W9576;
wire W9577;
wire W9578;
wire W9579;
wire W9580;
wire W9581;
wire W9582;
wire W9583;
wire W9584;
wire W9585;
wire W9586;
wire W9587;
wire W9588;
wire W9589;
wire W9590;
wire W9591;
wire W9592;
wire W9593;
wire W9594;
wire W9595;
wire W9596;
wire W9597;
wire W9598;
wire W9599;
wire W9600;
wire W9601;
wire W9602;
wire W9603;
wire W9604;
wire W9605;
wire W9606;
wire W9607;
wire W9608;
wire W9609;
wire W9610;
wire W9611;
wire W9612;
wire W9613;
wire W9614;
wire W9615;
wire W9616;
wire W9617;
wire W9618;
wire W9619;
wire W9620;
wire W9621;
wire W9622;
wire W9623;
wire W9624;
wire W9625;
wire W9626;
wire W9627;
wire W9628;
wire W9629;
wire W9630;
wire W9631;
wire W9632;
wire W9633;
wire W9634;
wire W9635;
wire W9636;
wire W9637;
wire W9638;
wire W9639;
wire W9640;
wire W9641;
wire W9642;
wire W9643;
wire W9644;
wire W9645;
wire W9646;
wire W9647;
wire W9648;
wire W9649;
wire W9650;
wire W9651;
wire W9652;
wire W9653;
wire W9654;
wire W9655;
wire W9656;
wire W9657;
wire W9658;
wire W9659;
wire W9660;
wire W9661;
wire W9662;
wire W9663;
wire W9664;
wire W9665;
wire W9666;
wire W9667;
wire W9668;
wire W9669;
wire W9670;
wire W9671;
wire W9672;
wire W9673;
wire W9674;
wire W9675;
wire W9676;
wire W9677;
wire W9678;
wire W9679;
wire W9680;
wire W9681;
wire W9682;
wire W9683;
wire W9684;
wire W9685;
wire W9686;
wire W9687;
wire W9688;
wire W9689;
wire W9690;
wire W9691;
wire W9692;
wire W9693;
wire W9694;
wire W9695;
wire W9696;
wire W9697;
wire W9698;
wire W9699;
wire W9700;
wire W9701;
wire W9702;
wire W9703;
wire W9704;
wire W9705;
wire W9706;
wire W9707;
wire W9708;
wire W9709;
wire W9710;
wire W9711;
wire W9712;
wire W9713;
wire W9714;
wire W9715;
wire W9716;
wire W9717;
wire W9718;
wire W9719;
wire W9720;
wire W9721;
wire W9722;
wire W9723;
wire W9724;
wire W9725;
wire W9726;
wire W9727;
wire W9728;
wire W9729;
wire W9730;
wire W9731;
wire W9732;
wire W9733;
wire W9734;
wire W9735;
wire W9736;
wire W9737;
wire W9738;
wire W9739;
wire W9740;
wire W9741;
wire W9742;
wire W9743;
wire W9744;
wire W9745;
wire W9746;
wire W9747;
wire W9748;
wire W9749;
wire W9750;
wire W9751;
wire W9752;
wire W9753;
wire W9754;
wire W9755;
wire W9756;
wire W9757;
wire W9758;
wire W9759;
wire W9760;
wire W9761;
wire W9762;
wire W9763;
wire W9764;
wire W9765;
wire W9766;
wire W9767;
wire W9768;
wire W9769;
wire W9770;
wire W9771;
wire W9772;
wire W9773;
wire W9774;
wire W9775;
wire W9776;
wire W9777;
wire W9778;
wire W9779;
wire W9780;
wire W9781;
wire W9782;
wire W9783;
wire W9784;
wire W9785;
wire W9786;
wire W9787;
wire W9788;
wire W9789;
wire W9790;
wire W9791;
wire W9792;
wire W9793;
wire W9794;
wire W9795;
wire W9796;
wire W9797;
wire W9798;
wire W9799;
wire W9800;
wire W9801;
wire W9802;
wire W9803;
wire W9804;
wire W9805;
wire W9806;
wire W9807;
wire W9808;
wire W9809;
wire W9810;
wire W9811;
wire W9812;
wire W9813;
wire W9814;
wire W9815;
wire W9816;
wire W9817;
wire W9818;
wire W9819;
wire W9820;
wire W9821;
wire W9822;
wire W9823;
wire W9824;
wire W9825;
wire W9826;
wire W9827;
wire W9828;
wire W9829;
wire W9830;
wire W9831;
wire W9832;
wire W9833;
wire W9834;
wire W9835;
wire W9836;
wire W9837;
wire W9838;
wire W9839;
wire W9840;
wire W9841;
wire W9842;
wire W9843;
wire W9844;
wire W9845;
wire W9846;
wire W9847;
wire W9848;
wire W9849;
wire W9850;
wire W9851;
wire W9852;
wire W9853;
wire W9854;
wire W9855;
wire W9856;
wire W9857;
wire W9858;
wire W9859;
wire W9860;
wire W9861;
wire W9862;
wire W9863;
wire W9864;
wire W9865;
wire W9866;
wire W9867;
wire W9868;
wire W9869;
wire W9870;
wire W9871;
wire W9872;
wire W9873;
wire W9874;
wire W9875;
wire W9876;
wire W9877;
wire W9878;
wire W9879;
wire W9880;
wire W9881;
wire W9882;
wire W9883;
wire W9884;
wire W9885;
wire W9886;
wire W9887;
wire W9888;
wire W9889;
wire W9890;
wire W9891;
wire W9892;
wire W9893;
wire W9894;
wire W9895;
wire W9896;
wire W9897;
wire W9898;
wire W9899;
wire W9900;
wire W9901;
wire W9902;
wire W9903;
wire W9904;
wire W9905;
wire W9906;
wire W9907;
wire W9908;
wire W9909;
wire W9910;
wire W9911;
wire W9912;
wire W9913;
wire W9914;
wire W9915;
wire W9916;
wire W9917;
wire W9918;
wire W9919;
wire W9920;
wire W9921;
wire W9922;
wire W9923;
wire W9924;
wire W9925;
wire W9926;
wire W9927;
wire W9928;
wire W9929;
wire W9930;
wire W9931;
wire W9932;
wire W9933;
wire W9934;
wire W9935;
wire W9936;
wire W9937;
wire W9938;
wire W9939;
wire W9940;
wire W9941;
wire W9942;
wire W9943;
wire W9944;
wire W9945;
wire W9946;
wire W9947;
wire W9948;
wire W9949;
wire W9950;
wire W9951;
wire W9952;
wire W9953;
wire W9954;
wire W9955;
wire W9956;
wire W9957;
wire W9958;
wire W9959;
wire W9960;
wire W9961;
wire W9962;
wire W9963;
wire W9964;
wire W9965;
wire W9966;
wire W9967;
wire W9968;
wire W9969;
wire W9970;
wire W9971;
wire W9972;
wire W9973;
wire W9974;
wire W9975;
wire W9976;
wire W9977;
wire W9978;
wire W9979;
wire W9980;
wire W9981;
wire W9982;
wire W9983;
wire W9984;
wire W9985;
wire W9986;
wire W9987;
wire W9988;
wire W9989;
wire W9990;
wire W9991;
wire W9992;
wire W9993;
wire W9994;
wire W9995;
wire W9996;
wire W9997;
wire W9998;
wire W9999;
wire W10000;
wire W10001;
wire W10002;
wire W10003;
wire W10004;
wire W10005;
wire W10006;
wire W10007;
wire W10008;
wire W10009;
wire W10010;
wire W10011;
wire W10012;
wire W10013;
wire W10014;
wire W10015;
wire W10016;
wire W10017;
wire W10018;
wire W10019;
wire W10020;
wire W10021;
wire W10022;
wire W10023;
wire W10024;
wire W10025;
wire W10026;
wire W10027;
wire W10028;
wire W10029;
wire W10030;
wire W10031;
wire W10032;
wire W10033;
wire W10034;
wire W10035;
wire W10036;
wire W10037;
wire W10038;
wire W10039;
wire W10040;
wire W10041;
wire W10042;
wire W10043;
wire W10044;
wire W10045;
wire W10046;
wire W10047;
wire W10048;
wire W10049;
wire W10050;
wire W10051;
wire W10052;
wire W10053;
wire W10054;
wire W10055;
wire W10056;
wire W10057;
wire W10058;
wire W10059;
wire W10060;
wire W10061;
wire W10062;
wire W10063;
wire W10064;
wire W10065;
wire W10066;
wire W10067;
wire W10068;
wire W10069;
wire W10070;
wire W10071;
wire W10072;
wire W10073;
wire W10074;
wire W10075;
wire W10076;
wire W10077;
wire W10078;
wire W10079;
wire W10080;
wire W10081;
wire W10082;
wire W10083;
wire W10084;
wire W10085;
wire W10086;
wire W10087;
wire W10088;
wire W10089;
wire W10090;
wire W10091;
wire W10092;
wire W10093;
wire W10094;
wire W10095;
wire W10096;
wire W10097;
wire W10098;
wire W10099;
wire W10100;
wire W10101;
wire W10102;
wire W10103;
wire W10104;
wire W10105;
wire W10106;
wire W10107;
wire W10108;
wire W10109;
wire W10110;
wire W10111;
wire W10112;
wire W10113;
wire W10114;
wire W10115;
wire W10116;
wire W10117;
wire W10118;
wire W10119;
wire W10120;
wire W10121;
wire W10122;
wire W10123;
wire W10124;
wire W10125;
wire W10126;
wire W10127;
wire W10128;
wire W10129;
wire W10130;
wire W10131;
wire W10132;
wire W10133;
wire W10134;
wire W10135;
wire W10136;
wire W10137;
wire W10138;
wire W10139;
wire W10140;
wire W10141;
wire W10142;
wire W10143;
wire W10144;
wire W10145;
wire W10146;
wire W10147;
wire W10148;
wire W10149;
wire W10150;
wire W10151;
wire W10152;
wire W10153;
wire W10154;
wire W10155;
wire W10156;
wire W10157;
wire W10158;
wire W10159;
wire W10160;
wire W10161;
wire W10162;
wire W10163;
wire W10164;
wire W10165;
wire W10166;
wire W10167;
wire W10168;
wire W10169;
wire W10170;
wire W10171;
wire W10172;
wire W10173;
wire W10174;
wire W10175;
wire W10176;
wire W10177;
wire W10178;
wire W10179;
wire W10180;
wire W10181;
wire W10182;
wire W10183;
wire W10184;
wire W10185;
wire W10186;
wire W10187;
wire W10188;
wire W10189;
wire W10190;
wire W10191;
wire W10192;
wire W10193;
wire W10194;
wire W10195;
wire W10196;
wire W10197;
wire W10198;
wire W10199;
wire W10200;
wire W10201;
wire W10202;
wire W10203;
wire W10204;
wire W10205;
wire W10206;
wire W10207;
wire W10208;
wire W10209;
wire W10210;
wire W10211;
wire W10212;
wire W10213;
wire W10214;
wire W10215;
wire W10216;
wire W10217;
wire W10218;
wire W10219;
wire W10220;
wire W10221;
wire W10222;
wire W10223;
wire W10224;
wire W10225;
wire W10226;
wire W10227;
wire W10228;
wire W10229;
wire W10230;
wire W10231;
wire W10232;
wire W10233;
wire W10234;
wire W10235;
wire W10236;
wire W10237;
wire W10238;
wire W10239;
wire W10240;
wire W10241;
wire W10242;
wire W10243;
wire W10244;
wire W10245;
wire W10246;
wire W10247;
wire W10248;
wire W10249;
wire W10250;
wire W10251;
wire W10252;
wire W10253;
wire W10254;
wire W10255;
wire W10256;
wire W10257;
wire W10258;
wire W10259;
wire W10260;
wire W10261;
wire W10262;
wire W10263;
wire W10264;
wire W10265;
wire W10266;
wire W10267;
wire W10268;
wire W10269;
wire W10270;
wire W10271;
wire W10272;
wire W10273;
wire W10274;
wire W10275;
wire W10276;
wire W10277;
wire W10278;
wire W10279;
wire W10280;
wire W10281;
wire W10282;
wire W10283;
wire W10284;
wire W10285;
wire W10286;
wire W10287;
wire W10288;
wire W10289;
wire W10290;
wire W10291;
wire W10292;
wire W10293;
wire W10294;
wire W10295;
wire W10296;
wire W10297;
wire W10298;
wire W10299;
wire W10300;
wire W10301;
wire W10302;
wire W10303;
wire W10304;
wire W10305;
wire W10306;
wire W10307;
wire W10308;
wire W10309;
wire W10310;
wire W10311;
wire W10312;
wire W10313;
wire W10314;
wire W10315;
wire W10316;
wire W10317;
wire W10318;
wire W10319;
wire W10320;
wire W10321;
wire W10322;
wire W10323;
wire W10324;
wire W10325;
wire W10326;
wire W10327;
wire W10328;
wire W10329;
wire W10330;
wire W10331;
wire W10332;
wire W10333;
wire W10334;
wire W10335;
wire W10336;
wire W10337;
wire W10338;
wire W10339;
wire W10340;
wire W10341;
wire W10342;
wire W10343;
wire W10344;
wire W10345;
wire W10346;
wire W10347;
wire W10348;
wire W10349;
wire W10350;
wire W10351;
wire W10352;
wire W10353;
wire W10354;
wire W10355;
wire W10356;
wire W10357;
wire W10358;
wire W10359;
wire W10360;
wire W10361;
wire W10362;
wire W10363;
wire W10364;
wire W10365;
wire W10366;
wire W10367;
wire W10368;
wire W10369;
wire W10370;
wire W10371;
wire W10372;
wire W10373;
wire W10374;
wire W10375;
wire W10376;
wire W10377;
wire W10378;
wire W10379;
wire W10380;
wire W10381;
wire W10382;
wire W10383;
wire W10384;
wire W10385;
wire W10386;
wire W10387;
wire W10388;
wire W10389;
wire W10390;
wire W10391;
wire W10392;
wire W10393;
wire W10394;
wire W10395;
wire W10396;
wire W10397;
wire W10398;
wire W10399;
wire W10400;
wire W10401;
wire W10402;
wire W10403;
wire W10404;
wire W10405;
wire W10406;
wire W10407;
wire W10408;
wire W10409;
wire W10410;
wire W10411;
wire W10412;
wire W10413;
wire W10414;
wire W10415;
wire W10416;
wire W10417;
wire W10418;
wire W10419;
wire W10420;
wire W10421;
wire W10422;
wire W10423;
wire W10424;
wire W10425;
wire W10426;
wire W10427;
wire W10428;
wire W10429;
wire W10430;
wire W10431;
wire W10432;
wire W10433;
wire W10434;
wire W10435;
wire W10436;
wire W10437;
wire W10438;
wire W10439;
wire W10440;
wire W10441;
wire W10442;
wire W10443;
wire W10444;
wire W10445;
wire W10446;
wire W10447;
wire W10448;
wire W10449;
wire W10450;
wire W10451;
wire W10452;
wire W10453;
wire W10454;
wire W10455;
wire W10456;
wire W10457;
wire W10458;
wire W10459;
wire W10460;
wire W10461;
wire W10462;
wire W10463;
wire W10464;
wire W10465;
wire W10466;
wire W10467;
wire W10468;
wire W10469;
wire W10470;
wire W10471;
wire W10472;
wire W10473;
wire W10474;
wire W10475;
wire W10476;
wire W10477;
wire W10478;
wire W10479;
wire W10480;
wire W10481;
wire W10482;
wire W10483;
wire W10484;
wire W10485;
wire W10486;
wire W10487;
wire W10488;
wire W10489;
wire W10490;
wire W10491;
wire W10492;
wire W10493;
wire W10494;
wire W10495;
wire W10496;
wire W10497;
wire W10498;
wire W10499;
wire W10500;
wire W10501;
wire W10502;
wire W10503;
wire W10504;
wire W10505;
wire W10506;
wire W10507;
wire W10508;
wire W10509;
wire W10510;
wire W10511;
wire W10512;
wire W10513;
wire W10514;
wire W10515;
wire W10516;
wire W10517;
wire W10518;
wire W10519;
wire W10520;
wire W10521;
wire W10522;
wire W10523;
wire W10524;
wire W10525;
wire W10526;
wire W10527;
wire W10528;
wire W10529;
wire W10530;
wire W10531;
wire W10532;
wire W10533;
wire W10534;
wire W10535;
wire W10536;
wire W10537;
wire W10538;
wire W10539;
wire W10540;
wire W10541;
wire W10542;
wire W10543;
wire W10544;
wire W10545;
wire W10546;
wire W10547;
wire W10548;
wire W10549;
wire W10550;
wire W10551;
wire W10552;
wire W10553;
wire W10554;
wire W10555;
wire W10556;
wire W10557;
wire W10558;
wire W10559;
wire W10560;
wire W10561;
wire W10562;
wire W10563;
wire W10564;
wire W10565;
wire W10566;
wire W10567;
wire W10568;
wire W10569;
wire W10570;
wire W10571;
wire W10572;
wire W10573;
wire W10574;
wire W10575;
wire W10576;
wire W10577;
wire W10578;
wire W10579;
wire W10580;
wire W10581;
wire W10582;
wire W10583;
wire W10584;
wire W10585;
wire W10586;
wire W10587;
wire W10588;
wire W10589;
wire W10590;
wire W10591;
wire W10592;
wire W10593;
wire W10594;
wire W10595;
wire W10596;
wire W10597;
wire W10598;
wire W10599;
wire W10600;
wire W10601;
wire W10602;
wire W10603;
wire W10604;
wire W10605;
wire W10606;
wire W10607;
wire W10608;
wire W10609;
wire W10610;
wire W10611;
wire W10612;
wire W10613;
wire W10614;
wire W10615;
wire W10616;
wire W10617;
wire W10618;
wire W10619;
wire W10620;
wire W10621;
wire W10622;
wire W10623;
wire W10624;
wire W10625;
wire W10626;
wire W10627;
wire W10628;
wire W10629;
wire W10630;
wire W10631;
wire W10632;
wire W10633;
wire W10634;
wire W10635;
wire W10636;
wire W10637;
wire W10638;
wire W10639;
wire W10640;
wire W10641;
wire W10642;
wire W10643;
wire W10644;
wire W10645;
wire W10646;
wire W10647;
wire W10648;
wire W10649;
wire W10650;
wire W10651;
wire W10652;
wire W10653;
wire W10654;
wire W10655;
wire W10656;
wire W10657;
wire W10658;
wire W10659;
wire W10660;
wire W10661;
wire W10662;
wire W10663;
wire W10664;
wire W10665;
wire W10666;
wire W10667;
wire W10668;
wire W10669;
wire W10670;
wire W10671;
wire W10672;
wire W10673;
wire W10674;
wire W10675;
wire W10676;
wire W10677;
wire W10678;
wire W10679;
wire W10680;
wire W10681;
wire W10682;
wire W10683;
wire W10684;
wire W10685;
wire W10686;
wire W10687;
wire W10688;
wire W10689;
wire W10690;
wire W10691;
wire W10692;
wire W10693;
wire W10694;
wire W10695;
wire W10696;
wire W10697;
wire W10698;
wire W10699;
wire W10700;
wire W10701;
wire W10702;
wire W10703;
wire W10704;
wire W10705;
wire W10706;
wire W10707;
wire W10708;
wire W10709;
wire W10710;
wire W10711;
wire W10712;
wire W10713;
wire W10714;
wire W10715;
wire W10716;
wire W10717;
wire W10718;
wire W10719;
wire W10720;
wire W10721;
wire W10722;
wire W10723;
wire W10724;
wire W10725;
wire W10726;
wire W10727;
wire W10728;
wire W10729;
wire W10730;
wire W10731;
wire W10732;
wire W10733;
wire W10734;
wire W10735;
wire W10736;
wire W10737;
wire W10738;
wire W10739;
wire W10740;
wire W10741;
wire W10742;
wire W10743;
wire W10744;
wire W10745;
wire W10746;
wire W10747;
wire W10748;
wire W10749;
wire W10750;
wire W10751;
wire W10752;
wire W10753;
wire W10754;
wire W10755;
wire W10756;
wire W10757;
wire W10758;
wire W10759;
wire W10760;
wire W10761;
wire W10762;
wire W10763;
wire W10764;
wire W10765;
wire W10766;
wire W10767;
wire W10768;
wire W10769;
wire W10770;
wire W10771;
wire W10772;
wire W10773;
wire W10774;
wire W10775;
wire W10776;
wire W10777;
wire W10778;
wire W10779;
wire W10780;
wire W10781;
wire W10782;
wire W10783;
wire W10784;
wire W10785;
wire W10786;
wire W10787;
wire W10788;
wire W10789;
wire W10790;
wire W10791;
wire W10792;
wire W10793;
wire W10794;
wire W10795;
wire W10796;
wire W10797;
wire W10798;
wire W10799;
wire W10800;
wire W10801;
wire W10802;
wire W10803;
wire W10804;
wire W10805;
wire W10806;
wire W10807;
wire W10808;
wire W10809;
wire W10810;
wire W10811;
wire W10812;
wire W10813;
wire W10814;
wire W10815;
wire W10816;
wire W10817;
wire W10818;
wire W10819;
wire W10820;
wire W10821;
wire W10822;
wire W10823;
wire W10824;
wire W10825;
wire W10826;
wire W10827;
wire W10828;
wire W10829;
wire W10830;
wire W10831;
wire W10832;
wire W10833;
wire W10834;
wire W10835;
wire W10836;
wire W10837;
wire W10838;
wire W10839;
wire W10840;
wire W10841;
wire W10842;
wire W10843;
wire W10844;
wire W10845;
wire W10846;
wire W10847;
wire W10848;
wire W10849;
wire W10850;
wire W10851;
wire W10852;
wire W10853;
wire W10854;
wire W10855;
wire W10856;
wire W10857;
wire W10858;
wire W10859;
wire W10860;
wire W10861;
wire W10862;
wire W10863;
wire W10864;
wire W10865;
wire W10866;
wire W10867;
wire W10868;
wire W10869;
wire W10870;
wire W10871;
wire W10872;
wire W10873;
wire W10874;
wire W10875;
wire W10876;
wire W10877;
wire W10878;
wire W10879;
wire W10880;
wire W10881;
wire W10882;
wire W10883;
wire W10884;
wire W10885;
wire W10886;
wire W10887;
wire W10888;
wire W10889;
wire W10890;
wire W10891;
wire W10892;
wire W10893;
wire W10894;
wire W10895;
wire W10896;
wire W10897;
wire W10898;
wire W10899;
wire W10900;
wire W10901;
wire W10902;
wire W10903;
wire W10904;
wire W10905;
wire W10906;
wire W10907;
wire W10908;
wire W10909;
wire W10910;
wire W10911;
wire W10912;
wire W10913;
wire W10914;
wire W10915;
wire W10916;
wire W10917;
wire W10918;
wire W10919;
wire W10920;
wire W10921;
wire W10922;
wire W10923;
wire W10924;
wire W10925;
wire W10926;
wire W10927;
wire W10928;
wire W10929;
wire W10930;
wire W10931;
wire W10932;
wire W10933;
wire W10934;
wire W10935;
wire W10936;
wire W10937;
wire W10938;
wire W10939;
wire W10940;
wire W10941;
wire W10942;
wire W10943;
wire W10944;
wire W10945;
wire W10946;
wire W10947;
wire W10948;
wire W10949;
wire W10950;
wire W10951;
wire W10952;
wire W10953;
wire W10954;
wire W10955;
wire W10956;
wire W10957;
wire W10958;
wire W10959;
wire W10960;
wire W10961;
wire W10962;
wire W10963;
wire W10964;
wire W10965;
wire W10966;
wire W10967;
wire W10968;
wire W10969;
wire W10970;
wire W10971;
wire W10972;
wire W10973;
wire W10974;
wire W10975;
wire W10976;
wire W10977;
wire W10978;
wire W10979;
wire W10980;
wire W10981;
wire W10982;
wire W10983;
wire W10984;
wire W10985;
wire W10986;
wire W10987;
wire W10988;
wire W10989;
wire W10990;
wire W10991;
wire W10992;
wire W10993;
wire W10994;
wire W10995;
wire W10996;
wire W10997;
wire W10998;
wire W10999;
wire W11000;
wire W11001;
wire W11002;
wire W11003;
wire W11004;
wire W11005;
wire W11006;
wire W11007;
wire W11008;
wire W11009;
wire W11010;
wire W11011;
wire W11012;
wire W11013;
wire W11014;
wire W11015;
wire W11016;
wire W11017;
wire W11018;
wire W11019;
wire W11020;
wire W11021;
wire W11022;
wire W11023;
wire W11024;
wire W11025;
wire W11026;
wire W11027;
wire W11028;
wire W11029;
wire W11030;
wire W11031;
wire W11032;
wire W11033;
wire W11034;
wire W11035;
wire W11036;
wire W11037;
wire W11038;
wire W11039;
wire W11040;
wire W11041;
wire W11042;
wire W11043;
wire W11044;
wire W11045;
wire W11046;
wire W11047;
wire W11048;
wire W11049;
wire W11050;
wire W11051;
wire W11052;
wire W11053;
wire W11054;
wire W11055;
wire W11056;
wire W11057;
wire W11058;
wire W11059;
wire W11060;
wire W11061;
wire W11062;
wire W11063;
wire W11064;
wire W11065;
wire W11066;
wire W11067;
wire W11068;
wire W11069;
wire W11070;
wire W11071;
wire W11072;
wire W11073;
wire W11074;
wire W11075;
wire W11076;
wire W11077;
wire W11078;
wire W11079;
wire W11080;
wire W11081;
wire W11082;
wire W11083;
wire W11084;
wire W11085;
wire W11086;
wire W11087;
wire W11088;
wire W11089;
wire W11090;
wire W11091;
wire W11092;
wire W11093;
wire W11094;
wire W11095;
wire W11096;
wire W11097;
wire W11098;
wire W11099;
wire W11100;
wire W11101;
wire W11102;
wire W11103;
wire W11104;
wire W11105;
wire W11106;
wire W11107;
wire W11108;
wire W11109;
wire W11110;
wire W11111;
wire W11112;
wire W11113;
wire W11114;
wire W11115;
wire W11116;
wire W11117;
wire W11118;
wire W11119;
wire W11120;
wire W11121;
wire W11122;
wire W11123;
wire W11124;
wire W11125;
wire W11126;
wire W11127;
wire W11128;
wire W11129;
wire W11130;
wire W11131;
wire W11132;
wire W11133;
wire W11134;
wire W11135;
wire W11136;
wire W11137;
wire W11138;
wire W11139;
wire W11140;
wire W11141;
wire W11142;
wire W11143;
wire W11144;
wire W11145;
wire W11146;
wire W11147;
wire W11148;
wire W11149;
wire W11150;
wire W11151;
wire W11152;
wire W11153;
wire W11154;
wire W11155;
wire W11156;
wire W11157;
wire W11158;
wire W11159;
wire W11160;
wire W11161;
wire W11162;
wire W11163;
wire W11164;
wire W11165;
wire W11166;
wire W11167;
wire W11168;
wire W11169;
wire W11170;
wire W11171;
wire W11172;
wire W11173;
wire W11174;
wire W11175;
wire W11176;
wire W11177;
wire W11178;
wire W11179;
wire W11180;
wire W11181;
wire W11182;
wire W11183;
wire W11184;
wire W11185;
wire W11186;
wire W11187;
wire W11188;
wire W11189;
wire W11190;
wire W11191;
wire W11192;
wire W11193;
wire W11194;
wire W11195;
wire W11196;
wire W11197;
wire W11198;
wire W11199;
wire W11200;
wire W11201;
wire W11202;
wire W11203;
wire W11204;
wire W11205;
wire W11206;
wire W11207;
wire W11208;
wire W11209;
wire W11210;
wire W11211;
wire W11212;
wire W11213;
wire W11214;
wire W11215;
wire W11216;
wire W11217;
wire W11218;
wire W11219;
wire W11220;
wire W11221;
wire W11222;
wire W11223;
wire W11224;
wire W11225;
wire W11226;
wire W11227;
wire W11228;
wire W11229;
wire W11230;
wire W11231;
wire W11232;
wire W11233;
wire W11234;
wire W11235;
wire W11236;
wire W11237;
wire W11238;
wire W11239;
wire W11240;
wire W11241;
wire W11242;
wire W11243;
wire W11244;
wire W11245;
wire W11246;
wire W11247;
wire W11248;
wire W11249;
wire W11250;
wire W11251;
wire W11252;
wire W11253;
wire W11254;
wire W11255;
wire W11256;
wire W11257;
wire W11258;
wire W11259;
wire W11260;
wire W11261;
wire W11262;
wire W11263;
wire W11264;
wire W11265;
wire W11266;
wire W11267;
wire W11268;
wire W11269;
wire W11270;
wire W11271;
wire W11272;
wire W11273;
wire W11274;
wire W11275;
wire W11276;
wire W11277;
wire W11278;
wire W11279;
wire W11280;
wire W11281;
wire W11282;
wire W11283;
wire W11284;
wire W11285;
wire W11286;
wire W11287;
wire W11288;
wire W11289;
wire W11290;
wire W11291;
wire W11292;
wire W11293;
wire W11294;
wire W11295;
wire W11296;
wire W11297;
wire W11298;
wire W11299;
wire W11300;
wire W11301;
wire W11302;
wire W11303;
wire W11304;
wire W11305;
wire W11306;
wire W11307;
wire W11308;
wire W11309;
wire W11310;
wire W11311;
wire W11312;
wire W11313;
wire W11314;
wire W11315;
wire W11316;
wire W11317;
wire W11318;
wire W11319;
wire W11320;
wire W11321;
wire W11322;
wire W11323;
wire W11324;
wire W11325;
wire W11326;
wire W11327;
wire W11328;
wire W11329;
wire W11330;
wire W11331;
wire W11332;
wire W11333;
wire W11334;
wire W11335;
wire W11336;
wire W11337;
wire W11338;
wire W11339;
wire W11340;
wire W11341;
wire W11342;
wire W11343;
wire W11344;
wire W11345;
wire W11346;
wire W11347;
wire W11348;
wire W11349;
wire W11350;
wire W11351;
wire W11352;
wire W11353;
wire W11354;
wire W11355;
wire W11356;
wire W11357;
wire W11358;
wire W11359;
wire W11360;
wire W11361;
wire W11362;
wire W11363;
wire W11364;
wire W11365;
wire W11366;
wire W11367;
wire W11368;
wire W11369;
wire W11370;
wire W11371;
wire W11372;
wire W11373;
wire W11374;
wire W11375;
wire W11376;
wire W11377;
wire W11378;
wire W11379;
wire W11380;
wire W11381;
wire W11382;
wire W11383;
wire W11384;
wire W11385;
wire W11386;
wire W11387;
wire W11388;
wire W11389;
wire W11390;
wire W11391;
wire W11392;
wire W11393;
wire W11394;
wire W11395;
wire W11396;
wire W11397;
wire W11398;
wire W11399;
wire W11400;
wire W11401;
wire W11402;
wire W11403;
wire W11404;
wire W11405;
wire W11406;
wire W11407;
wire W11408;
wire W11409;
wire W11410;
wire W11411;
wire W11412;
wire W11413;
wire W11414;
wire W11415;
wire W11416;
wire W11417;
wire W11418;
wire W11419;
wire W11420;
wire W11421;
wire W11422;
wire W11423;
wire W11424;
wire W11425;
wire W11426;
wire W11427;
wire W11428;
wire W11429;
wire W11430;
wire W11431;
wire W11432;
wire W11433;
wire W11434;
wire W11435;
wire W11436;
wire W11437;
wire W11438;
wire W11439;
wire W11440;
wire W11441;
wire W11442;
wire W11443;
wire W11444;
wire W11445;
wire W11446;
wire W11447;
wire W11448;
wire W11449;
wire W11450;
wire W11451;
wire W11452;
wire W11453;
wire W11454;
wire W11455;
wire W11456;
wire W11457;
wire W11458;
wire W11459;
wire W11460;
wire W11461;
wire W11462;
wire W11463;
wire W11464;
wire W11465;
wire W11466;
wire W11467;
wire W11468;
wire W11469;
wire W11470;
wire W11471;
wire W11472;
wire W11473;
wire W11474;
wire W11475;
wire W11476;
wire W11477;
wire W11478;
wire W11479;
wire W11480;
wire W11481;
wire W11482;
wire W11483;
wire W11484;
wire W11485;
wire W11486;
wire W11487;
wire W11488;
wire W11489;
wire W11490;
wire W11491;
wire W11492;
wire W11493;
wire W11494;
wire W11495;
wire W11496;
wire W11497;
wire W11498;
wire W11499;
wire W11500;
wire W11501;
wire W11502;
wire W11503;
wire W11504;
wire W11505;
wire W11506;
wire W11507;
wire W11508;
wire W11509;
wire W11510;
wire W11511;
wire W11512;
wire W11513;
wire W11514;
wire W11515;
wire W11516;
wire W11517;
wire W11518;
wire W11519;
wire W11520;
wire W11521;
wire W11522;
wire W11523;
wire W11524;
wire W11525;
wire W11526;
wire W11527;
wire W11528;
wire W11529;
wire W11530;
wire W11531;
wire W11532;
wire W11533;
wire W11534;
wire W11535;
wire W11536;
wire W11537;
wire W11538;
wire W11539;
wire W11540;
wire W11541;
wire W11542;
wire W11543;
wire W11544;
wire W11545;
wire W11546;
wire W11547;
wire W11548;
wire W11549;
wire W11550;
wire W11551;
wire W11552;
wire W11553;
wire W11554;
wire W11555;
wire W11556;
wire W11557;
wire W11558;
wire W11559;
wire W11560;
wire W11561;
wire W11562;
wire W11563;
wire W11564;
wire W11565;
wire W11566;
wire W11567;
wire W11568;
wire W11569;
wire W11570;
wire W11571;
wire W11572;
wire W11573;
wire W11574;
wire W11575;
wire W11576;
wire W11577;
wire W11578;
wire W11579;
wire W11580;
wire W11581;
wire W11582;
wire W11583;
wire W11584;
wire W11585;
wire W11586;
wire W11587;
wire W11588;
wire W11589;
wire W11590;
wire W11591;
wire W11592;
wire W11593;
wire W11594;
wire W11595;
wire W11596;
wire W11597;
wire W11598;
wire W11599;
wire W11600;
wire W11601;
wire W11602;
wire W11603;
wire W11604;
wire W11605;
wire W11606;
wire W11607;
wire W11608;
wire W11609;
wire W11610;
wire W11611;
wire W11612;
wire W11613;
wire W11614;
wire W11615;
wire W11616;
wire W11617;
wire W11618;
wire W11619;
wire W11620;
wire W11621;
wire W11622;
wire W11623;
wire W11624;
wire W11625;
wire W11626;
wire W11627;
wire W11628;
wire W11629;
wire W11630;
wire W11631;
wire W11632;
wire W11633;
wire W11634;
wire W11635;
wire W11636;
wire W11637;
wire W11638;
wire W11639;
wire W11640;
wire W11641;
wire W11642;
wire W11643;
wire W11644;
wire W11645;
wire W11646;
wire W11647;
wire W11648;
wire W11649;
wire W11650;
wire W11651;
wire W11652;
wire W11653;
wire W11654;
wire W11655;
wire W11656;
wire W11657;
wire W11658;
wire W11659;
wire W11660;
wire W11661;
wire W11662;
wire W11663;
wire W11664;
wire W11665;
wire W11666;
wire W11667;
wire W11668;
wire W11669;
wire W11670;
wire W11671;
wire W11672;
wire W11673;
wire W11674;
wire W11675;
wire W11676;
wire W11677;
wire W11678;
wire W11679;
wire W11680;
wire W11681;
wire W11682;
wire W11683;
wire W11684;
wire W11685;
wire W11686;
wire W11687;
wire W11688;
wire W11689;
wire W11690;
wire W11691;
wire W11692;
wire W11693;
wire W11694;
wire W11695;
wire W11696;
wire W11697;
wire W11698;
wire W11699;
wire W11700;
wire W11701;
wire W11702;
wire W11703;
wire W11704;
wire W11705;
wire W11706;
wire W11707;
wire W11708;
wire W11709;
wire W11710;
wire W11711;
wire W11712;
wire W11713;
wire W11714;
wire W11715;
wire W11716;
wire W11717;
wire W11718;
wire W11719;
wire W11720;
wire W11721;
wire W11722;
wire W11723;
wire W11724;
wire W11725;
wire W11726;
wire W11727;
wire W11728;
wire W11729;
wire W11730;
wire W11731;
wire W11732;
wire W11733;
wire W11734;
wire W11735;
wire W11736;
wire W11737;
wire W11738;
wire W11739;
wire W11740;
wire W11741;
wire W11742;
wire W11743;
wire W11744;
wire W11745;
wire W11746;
wire W11747;
wire W11748;
wire W11749;
wire W11750;
wire W11751;
wire W11752;
wire W11753;
wire W11754;
wire W11755;
wire W11756;
wire W11757;
wire W11758;
wire W11759;
wire W11760;
wire W11761;
wire W11762;
wire W11763;
wire W11764;
wire W11765;
wire W11766;
wire W11767;
wire W11768;
wire W11769;
wire W11770;
wire W11771;
wire W11772;
wire W11773;
wire W11774;
wire W11775;
wire W11776;
wire W11777;
wire W11778;
wire W11779;
wire W11780;
wire W11781;
wire W11782;
wire W11783;
wire W11784;
wire W11785;
wire W11786;
wire W11787;
wire W11788;
wire W11789;
wire W11790;
wire W11791;
wire W11792;
wire W11793;
wire W11794;
wire W11795;
wire W11796;
wire W11797;
wire W11798;
wire W11799;
wire W11800;
wire W11801;
wire W11802;
wire W11803;
wire W11804;
wire W11805;
wire W11806;
wire W11807;
wire W11808;
wire W11809;
wire W11810;
wire W11811;
wire W11812;
wire W11813;
wire W11814;
wire W11815;
wire W11816;
wire W11817;
wire W11818;
wire W11819;
wire W11820;
wire W11821;
wire W11822;
wire W11823;
wire W11824;
wire W11825;
wire W11826;
wire W11827;
wire W11828;
wire W11829;
wire W11830;
wire W11831;
wire W11832;
wire W11833;
wire W11834;
wire W11835;
wire W11836;
wire W11837;
wire W11838;
wire W11839;
wire W11840;
wire W11841;
wire W11842;
wire W11843;
wire W11844;
wire W11845;
wire W11846;
wire W11847;
wire W11848;
wire W11849;
wire W11850;
wire W11851;
wire W11852;
wire W11853;
wire W11854;
wire W11855;
wire W11856;
wire W11857;
wire W11858;
wire W11859;
wire W11860;
wire W11861;
wire W11862;
wire W11863;
wire W11864;
wire W11865;
wire W11866;
wire W11867;
wire W11868;
wire W11869;
wire W11870;
wire W11871;
wire W11872;
wire W11873;
wire W11874;
wire W11875;
wire W11876;
wire W11877;
wire W11878;
wire W11879;
wire W11880;
wire W11881;
wire W11882;
wire W11883;
wire W11884;
wire W11885;
wire W11886;
wire W11887;
wire W11888;
wire W11889;
wire W11890;
wire W11891;
wire W11892;
wire W11893;
wire W11894;
wire W11895;
wire W11896;
wire W11897;
wire W11898;
wire W11899;
wire W11900;
wire W11901;
wire W11902;
wire W11903;
wire W11904;
wire W11905;
wire W11906;
wire W11907;
wire W11908;
wire W11909;
wire W11910;
wire W11911;
wire W11912;
wire W11913;
wire W11914;
wire W11915;
wire W11916;
wire W11917;
wire W11918;
wire W11919;
wire W11920;
wire W11921;
wire W11922;
wire W11923;
wire W11924;
wire W11925;
wire W11926;
wire W11927;
wire W11928;
wire W11929;
wire W11930;
wire W11931;
wire W11932;
wire W11933;
wire W11934;
wire W11935;
wire W11936;
wire W11937;
wire W11938;
wire W11939;
wire W11940;
wire W11941;
wire W11942;
wire W11943;
wire W11944;
wire W11945;
wire W11946;
wire W11947;
wire W11948;
wire W11949;
wire W11950;
wire W11951;
wire W11952;
wire W11953;
wire W11954;
wire W11955;
wire W11956;
wire W11957;
wire W11958;
wire W11959;
wire W11960;
wire W11961;
wire W11962;
wire W11963;
wire W11964;
wire W11965;
wire W11966;
wire W11967;
wire W11968;
wire W11969;
wire W11970;
wire W11971;
wire W11972;
wire W11973;
wire W11974;
wire W11975;
wire W11976;
wire W11977;
wire W11978;
wire W11979;
wire W11980;
wire W11981;
wire W11982;
wire W11983;
wire W11984;
wire W11985;
wire W11986;
wire W11987;
wire W11988;
wire W11989;
wire W11990;
wire W11991;
wire W11992;
wire W11993;
wire W11994;
wire W11995;
wire W11996;
wire W11997;
wire W11998;
wire W11999;
wire W12000;
wire W12001;
wire W12002;
wire W12003;
wire W12004;
wire W12005;
wire W12006;
wire W12007;
wire W12008;
wire W12009;
wire W12010;
wire W12011;
wire W12012;
wire W12013;
wire W12014;
wire W12015;
wire W12016;
wire W12017;
wire W12018;
wire W12019;
wire W12020;
wire W12021;
wire W12022;
wire W12023;
wire W12024;
wire W12025;
wire W12026;
wire W12027;
wire W12028;
wire W12029;
wire W12030;
wire W12031;
wire W12032;
wire W12033;
wire W12034;
wire W12035;
wire W12036;
wire W12037;
wire W12038;
wire W12039;
wire W12040;
wire W12041;
wire W12042;
wire W12043;
wire W12044;
wire W12045;
wire W12046;
wire W12047;
wire W12048;
wire W12049;
wire W12050;
wire W12051;
wire W12052;
wire W12053;
wire W12054;
wire W12055;
wire W12056;
wire W12057;
wire W12058;
wire W12059;
wire W12060;
wire W12061;
wire W12062;
wire W12063;
wire W12064;
wire W12065;
wire W12066;
wire W12067;
wire W12068;
wire W12069;
wire W12070;
wire W12071;
wire W12072;
wire W12073;
wire W12074;
wire W12075;
wire W12076;
wire W12077;
wire W12078;
wire W12079;
wire W12080;
wire W12081;
wire W12082;
wire W12083;
wire W12084;
wire W12085;
wire W12086;
wire W12087;
wire W12088;
wire W12089;
wire W12090;
wire W12091;
wire W12092;
wire W12093;
wire W12094;
wire W12095;
wire W12096;
wire W12097;
wire W12098;
wire W12099;
wire W12100;
wire W12101;
wire W12102;
wire W12103;
wire W12104;
wire W12105;
wire W12106;
wire W12107;
wire W12108;
wire W12109;
wire W12110;
wire W12111;
wire W12112;
wire W12113;
wire W12114;
wire W12115;
wire W12116;
wire W12117;
wire W12118;
wire W12119;
wire W12120;
wire W12121;
wire W12122;
wire W12123;
wire W12124;
wire W12125;
wire W12126;
wire W12127;
wire W12128;
wire W12129;
wire W12130;
wire W12131;
wire W12132;
wire W12133;
wire W12134;
wire W12135;
wire W12136;
wire W12137;
wire W12138;
wire W12139;
wire W12140;
wire W12141;
wire W12142;
wire W12143;
wire W12144;
wire W12145;
wire W12146;
wire W12147;
wire W12148;
wire W12149;
wire W12150;
wire W12151;
wire W12152;
wire W12153;
wire W12154;
wire W12155;
wire W12156;
wire W12157;
wire W12158;
wire W12159;
wire W12160;
wire W12161;
wire W12162;
wire W12163;
wire W12164;
wire W12165;
wire W12166;
wire W12167;
wire W12168;
wire W12169;
wire W12170;
wire W12171;
wire W12172;
wire W12173;
wire W12174;
wire W12175;
wire W12176;
wire W12177;
wire W12178;
wire W12179;
wire W12180;
wire W12181;
wire W12182;
wire W12183;
wire W12184;
wire W12185;
wire W12186;
wire W12187;
wire W12188;
wire W12189;
wire W12190;
wire W12191;
wire W12192;
wire W12193;
wire W12194;
wire W12195;
wire W12196;
wire W12197;
wire W12198;
wire W12199;
wire W12200;
wire W12201;
wire W12202;
wire W12203;
wire W12204;
wire W12205;
wire W12206;
wire W12207;
wire W12208;
wire W12209;
wire W12210;
wire W12211;
wire W12212;
wire W12213;
wire W12214;
wire W12215;
wire W12216;
wire W12217;
wire W12218;
wire W12219;
wire W12220;
wire W12221;
wire W12222;
wire W12223;
wire W12224;
wire W12225;
wire W12226;
wire W12227;
wire W12228;
wire W12229;
wire W12230;
wire W12231;
wire W12232;
wire W12233;
wire W12234;
wire W12235;
wire W12236;
wire W12237;
wire W12238;
wire W12239;
wire W12240;
wire W12241;
wire W12242;
wire W12243;
wire W12244;
wire W12245;
wire W12246;
wire W12247;
wire W12248;
wire W12249;
wire W12250;
wire W12251;
wire W12252;
wire W12253;
wire W12254;
wire W12255;
wire W12256;
wire W12257;
wire W12258;
wire W12259;
wire W12260;
wire W12261;
wire W12262;
wire W12263;
wire W12264;
wire W12265;
wire W12266;
wire W12267;
wire W12268;
wire W12269;
wire W12270;
wire W12271;
wire W12272;
wire W12273;
wire W12274;
wire W12275;
wire W12276;
wire W12277;
wire W12278;
wire W12279;
wire W12280;
wire W12281;
wire W12282;
wire W12283;
wire W12284;
wire W12285;
wire W12286;
wire W12287;
wire W12288;
wire W12289;
wire W12290;
wire W12291;
wire W12292;
wire W12293;
wire W12294;
wire W12295;
wire W12296;
wire W12297;
wire W12298;
wire W12299;
wire W12300;
wire W12301;
wire W12302;
wire W12303;
wire W12304;
wire W12305;
wire W12306;
wire W12307;
wire W12308;
wire W12309;
wire W12310;
wire W12311;
wire W12312;
wire W12313;
wire W12314;
wire W12315;
wire W12316;
wire W12317;
wire W12318;
wire W12319;
wire W12320;
wire W12321;
wire W12322;
wire W12323;
wire W12324;
wire W12325;
wire W12326;
wire W12327;
wire W12328;
wire W12329;
wire W12330;
wire W12331;
wire W12332;
wire W12333;
wire W12334;
wire W12335;
wire W12336;
wire W12337;
wire W12338;
wire W12339;
wire W12340;
wire W12341;
wire W12342;
wire W12343;
wire W12344;
wire W12345;
wire W12346;
wire W12347;
wire W12348;
wire W12349;
wire W12350;
wire W12351;
wire W12352;
wire W12353;
wire W12354;
wire W12355;
wire W12356;
wire W12357;
wire W12358;
wire W12359;
wire W12360;
wire W12361;
wire W12362;
wire W12363;
wire W12364;
wire W12365;
wire W12366;
wire W12367;
wire W12368;
wire W12369;
wire W12370;
wire W12371;
wire W12372;
wire W12373;
wire W12374;
wire W12375;
wire W12376;
wire W12377;
wire W12378;
wire W12379;
wire W12380;
wire W12381;
wire W12382;
wire W12383;
wire W12384;
wire W12385;
wire W12386;
wire W12387;
wire W12388;
wire W12389;
wire W12390;
wire W12391;
wire W12392;
wire W12393;
wire W12394;
wire W12395;
wire W12396;
wire W12397;
wire W12398;
wire W12399;
wire W12400;
wire W12401;
wire W12402;
wire W12403;
wire W12404;
wire W12405;
wire W12406;
wire W12407;
wire W12408;
wire W12409;
wire W12410;
wire W12411;
wire W12412;
wire W12413;
wire W12414;
wire W12415;
wire W12416;
wire W12417;
wire W12418;
wire W12419;
wire W12420;
wire W12421;
wire W12422;
wire W12423;
wire W12424;
wire W12425;
wire W12426;
wire W12427;
wire W12428;
wire W12429;
wire W12430;
wire W12431;
wire W12432;
wire W12433;
wire W12434;
wire W12435;
wire W12436;
wire W12437;
wire W12438;
wire W12439;
wire W12440;
wire W12441;
wire W12442;
wire W12443;
wire W12444;
wire W12445;
wire W12446;
wire W12447;
wire W12448;
wire W12449;
wire W12450;
wire W12451;
wire W12452;
wire W12453;
wire W12454;
wire W12455;
wire W12456;
wire W12457;
wire W12458;
wire W12459;
wire W12460;
wire W12461;
wire W12462;
wire W12463;
wire W12464;
wire W12465;
wire W12466;
wire W12467;
wire W12468;
wire W12469;
wire W12470;
wire W12471;
wire W12472;
wire W12473;
wire W12474;
wire W12475;
wire W12476;
wire W12477;
wire W12478;
wire W12479;
wire W12480;
wire W12481;
wire W12482;
wire W12483;
wire W12484;
wire W12485;
wire W12486;
wire W12487;
wire W12488;
wire W12489;
wire W12490;
wire W12491;
wire W12492;
wire W12493;
wire W12494;
wire W12495;
wire W12496;
wire W12497;
wire W12498;
wire W12499;
wire W12500;
wire W12501;
wire W12502;
wire W12503;
wire W12504;
wire W12505;
wire W12506;
wire W12507;
wire W12508;
wire W12509;
wire W12510;
wire W12511;
wire W12512;
wire W12513;
wire W12514;
wire W12515;
wire W12516;
wire W12517;
wire W12518;
wire W12519;
wire W12520;
wire W12521;
wire W12522;
wire W12523;
wire W12524;
wire W12525;
wire W12526;
wire W12527;
wire W12528;
wire W12529;
wire W12530;
wire W12531;
wire W12532;
wire W12533;
wire W12534;
wire W12535;
wire W12536;
wire W12537;
wire W12538;
wire W12539;
wire W12540;
wire W12541;
wire W12542;
wire W12543;
wire W12544;
wire W12545;
wire W12546;
wire W12547;
wire W12548;
wire W12549;
wire W12550;
wire W12551;
wire W12552;
wire W12553;
wire W12554;
wire W12555;
wire W12556;
wire W12557;
wire W12558;
wire W12559;
wire W12560;
wire W12561;
wire W12562;
wire W12563;
wire W12564;
wire W12565;
wire W12566;
wire W12567;
wire W12568;
wire W12569;
wire W12570;
wire W12571;
wire W12572;
wire W12573;
wire W12574;
wire W12575;
wire W12576;
wire W12577;
wire W12578;
wire W12579;
wire W12580;
wire W12581;
wire W12582;
wire W12583;
wire W12584;
wire W12585;
wire W12586;
wire W12587;
wire W12588;
wire W12589;
wire W12590;
wire W12591;
wire W12592;
wire W12593;
wire W12594;
wire W12595;
wire W12596;
wire W12597;
wire W12598;
wire W12599;
wire W12600;
wire W12601;
wire W12602;
wire W12603;
wire W12604;
wire W12605;
wire W12606;
wire W12607;
wire W12608;
wire W12609;
wire W12610;
wire W12611;
wire W12612;
wire W12613;
wire W12614;
wire W12615;
wire W12616;
wire W12617;
wire W12618;
wire W12619;
wire W12620;
wire W12621;
wire W12622;
wire W12623;
wire W12624;
wire W12625;
wire W12626;
wire W12627;
wire W12628;
wire W12629;
wire W12630;
wire W12631;
wire W12632;
wire W12633;
wire W12634;
wire W12635;
wire W12636;
wire W12637;
wire W12638;
wire W12639;
wire W12640;
wire W12641;
wire W12642;
wire W12643;
wire W12644;
wire W12645;
wire W12646;
wire W12647;
wire W12648;
wire W12649;
wire W12650;
wire W12651;
wire W12652;
wire W12653;
wire W12654;
wire W12655;
wire W12656;
wire W12657;
wire W12658;
wire W12659;
wire W12660;
wire W12661;
wire W12662;
wire W12663;
wire W12664;
wire W12665;
wire W12666;
wire W12667;
wire W12668;
wire W12669;
wire W12670;
wire W12671;
wire W12672;
wire W12673;
wire W12674;
wire W12675;
wire W12676;
wire W12677;
wire W12678;
wire W12679;
wire W12680;
wire W12681;
wire W12682;
wire W12683;
wire W12684;
wire W12685;
wire W12686;
wire W12687;
wire W12688;
wire W12689;
wire W12690;
wire W12691;
wire W12692;
wire W12693;
wire W12694;
wire W12695;
wire W12696;
wire W12697;
wire W12698;
wire W12699;
wire W12700;
wire W12701;
wire W12702;
wire W12703;
wire W12704;
wire W12705;
wire W12706;
wire W12707;
wire W12708;
wire W12709;
wire W12710;
wire W12711;
wire W12712;
wire W12713;
wire W12714;
wire W12715;
wire W12716;
wire W12717;
wire W12718;
wire W12719;
wire W12720;
wire W12721;
wire W12722;
wire W12723;
wire W12724;
wire W12725;
wire W12726;
wire W12727;
wire W12728;
wire W12729;
wire W12730;
wire W12731;
wire W12732;
wire W12733;
wire W12734;
wire W12735;
wire W12736;
wire W12737;
wire W12738;
wire W12739;
wire W12740;
wire W12741;
wire W12742;
wire W12743;
wire W12744;
wire W12745;
wire W12746;
wire W12747;
wire W12748;
wire W12749;
wire W12750;
wire W12751;
wire W12752;
wire W12753;
wire W12754;
wire W12755;
wire W12756;
wire W12757;
wire W12758;
wire W12759;
wire W12760;
wire W12761;
wire W12762;
wire W12763;
wire W12764;
wire W12765;
wire W12766;
wire W12767;
wire W12768;
wire W12769;
wire W12770;
wire W12771;
wire W12772;
wire W12773;
wire W12774;
wire W12775;
wire W12776;
wire W12777;
wire W12778;
wire W12779;
wire W12780;
wire W12781;
wire W12782;
wire W12783;
wire W12784;
wire W12785;
wire W12786;
wire W12787;
wire W12788;
wire W12789;
wire W12790;
wire W12791;
wire W12792;
wire W12793;
wire W12794;
wire W12795;
wire W12796;
wire W12797;
wire W12798;
wire W12799;
wire W12800;
wire W12801;
wire W12802;
wire W12803;
wire W12804;
wire W12805;
wire W12806;
wire W12807;
wire W12808;
wire W12809;
wire W12810;
wire W12811;
wire W12812;
wire W12813;
wire W12814;
wire W12815;
wire W12816;
wire W12817;
wire W12818;
wire W12819;
wire W12820;
wire W12821;
wire W12822;
wire W12823;
wire W12824;
wire W12825;
wire W12826;
wire W12827;
wire W12828;
wire W12829;
wire W12830;
wire W12831;
wire W12832;
wire W12833;
wire W12834;
wire W12835;
wire W12836;
wire W12837;
wire W12838;
wire W12839;
wire W12840;
wire W12841;
wire W12842;
wire W12843;
wire W12844;
wire W12845;
wire W12846;
wire W12847;
wire W12848;
wire W12849;
wire W12850;
wire W12851;
wire W12852;
wire W12853;
wire W12854;
wire W12855;
wire W12856;
wire W12857;
wire W12858;
wire W12859;
wire W12860;
wire W12861;
wire W12862;
wire W12863;
wire W12864;
wire W12865;
wire W12866;
wire W12867;
wire W12868;
wire W12869;
wire W12870;
wire W12871;
wire W12872;
wire W12873;
wire W12874;
wire W12875;
wire W12876;
wire W12877;
wire W12878;
wire W12879;
wire W12880;
wire W12881;
wire W12882;
wire W12883;
wire W12884;
wire W12885;
wire W12886;
wire W12887;
wire W12888;
wire W12889;
wire W12890;
wire W12891;
wire W12892;
wire W12893;
wire W12894;
wire W12895;
wire W12896;
wire W12897;
wire W12898;
wire W12899;
wire W12900;
wire W12901;
wire W12902;
wire W12903;
wire W12904;
wire W12905;
wire W12906;
wire W12907;
wire W12908;
wire W12909;
wire W12910;
wire W12911;
wire W12912;
wire W12913;
wire W12914;
wire W12915;
wire W12916;
wire W12917;
wire W12918;
wire W12919;
wire W12920;
wire W12921;
wire W12922;
wire W12923;
wire W12924;
wire W12925;
wire W12926;
wire W12927;
wire W12928;
wire W12929;
wire W12930;
wire W12931;
wire W12932;
wire W12933;
wire W12934;
wire W12935;
wire W12936;
wire W12937;
wire W12938;
wire W12939;
wire W12940;
wire W12941;
wire W12942;
wire W12943;
wire W12944;
wire W12945;
wire W12946;
wire W12947;
wire W12948;
wire W12949;
wire W12950;
wire W12951;
wire W12952;
wire W12953;
wire W12954;
wire W12955;
wire W12956;
wire W12957;
wire W12958;
wire W12959;
wire W12960;
wire W12961;
wire W12962;
wire W12963;
wire W12964;
wire W12965;
wire W12966;
wire W12967;
wire W12968;
wire W12969;
wire W12970;
wire W12971;
wire W12972;
wire W12973;
wire W12974;
wire W12975;
wire W12976;
wire W12977;
wire W12978;
wire W12979;
wire W12980;
wire W12981;
wire W12982;
wire W12983;
wire W12984;
wire W12985;
wire W12986;
wire W12987;
wire W12988;
wire W12989;
wire W12990;
wire W12991;
wire W12992;
wire W12993;
wire W12994;
wire W12995;
wire W12996;
wire W12997;
wire W12998;
wire W12999;
wire W13000;
wire W13001;
wire W13002;
wire W13003;
wire W13004;
wire W13005;
wire W13006;
wire W13007;
wire W13008;
wire W13009;
wire W13010;
wire W13011;
wire W13012;
wire W13013;
wire W13014;
wire W13015;
wire W13016;
wire W13017;
wire W13018;
wire W13019;
wire W13020;
wire W13021;
wire W13022;
wire W13023;
wire W13024;
wire W13025;
wire W13026;
wire W13027;
wire W13028;
wire W13029;
wire W13030;
wire W13031;
wire W13032;
wire W13033;
wire W13034;
wire W13035;
wire W13036;
wire W13037;
wire W13038;
wire W13039;
wire W13040;
wire W13041;
wire W13042;
wire W13043;
wire W13044;
wire W13045;
wire W13046;
wire W13047;
wire W13048;
wire W13049;
wire W13050;
wire W13051;
wire W13052;
wire W13053;
wire W13054;
wire W13055;
wire W13056;
wire W13057;
wire W13058;
wire W13059;
wire W13060;
wire W13061;
wire W13062;
wire W13063;
wire W13064;
wire W13065;
wire W13066;
wire W13067;
wire W13068;
wire W13069;
wire W13070;
wire W13071;
wire W13072;
wire W13073;
wire W13074;
wire W13075;
wire W13076;
wire W13077;
wire W13078;
wire W13079;
wire W13080;
wire W13081;
wire W13082;
wire W13083;
wire W13084;
wire W13085;
wire W13086;
wire W13087;
wire W13088;
wire W13089;
wire W13090;
wire W13091;
wire W13092;
wire W13093;
wire W13094;
wire W13095;
wire W13096;
wire W13097;
wire W13098;
wire W13099;
wire W13100;
wire W13101;
wire W13102;
wire W13103;
wire W13104;
wire W13105;
wire W13106;
wire W13107;
wire W13108;
wire W13109;
wire W13110;
wire W13111;
wire W13112;
wire W13113;
wire W13114;
wire W13115;
wire W13116;
wire W13117;
wire W13118;
wire W13119;
wire W13120;
wire W13121;
wire W13122;
wire W13123;
wire W13124;
wire W13125;
wire W13126;
wire W13127;
wire W13128;
wire W13129;
wire W13130;
wire W13131;
wire W13132;
wire W13133;
wire W13134;
wire W13135;
wire W13136;
wire W13137;
wire W13138;
wire W13139;
wire W13140;
wire W13141;
wire W13142;
wire W13143;
wire W13144;
wire W13145;
wire W13146;
wire W13147;
wire W13148;
wire W13149;
wire W13150;
wire W13151;
wire W13152;
wire W13153;
wire W13154;
wire W13155;
wire W13156;
wire W13157;
wire W13158;
wire W13159;
wire W13160;
wire W13161;
wire W13162;
wire W13163;
wire W13164;
wire W13165;
wire W13166;
wire W13167;
wire W13168;
wire W13169;
wire W13170;
wire W13171;
wire W13172;
wire W13173;
wire W13174;
wire W13175;
wire W13176;
wire W13177;
wire W13178;
wire W13179;
wire W13180;
wire W13181;
wire W13182;
wire W13183;
wire W13184;
wire W13185;
wire W13186;
wire W13187;
wire W13188;
wire W13189;
wire W13190;
wire W13191;
wire W13192;
wire W13193;
wire W13194;
wire W13195;
wire W13196;
wire W13197;
wire W13198;
wire W13199;
wire W13200;
wire W13201;
wire W13202;
wire W13203;
wire W13204;
wire W13205;
wire W13206;
wire W13207;
wire W13208;
wire W13209;
wire W13210;
wire W13211;
wire W13212;
wire W13213;
wire W13214;
wire W13215;
wire W13216;
wire W13217;
wire W13218;
wire W13219;
wire W13220;
wire W13221;
wire W13222;
wire W13223;
wire W13224;
wire W13225;
wire W13226;
wire W13227;
wire W13228;
wire W13229;
wire W13230;
wire W13231;
wire W13232;
wire W13233;
wire W13234;
wire W13235;
wire W13236;
wire W13237;
wire W13238;
wire W13239;
wire W13240;
wire W13241;
wire W13242;
wire W13243;
wire W13244;
wire W13245;
wire W13246;
wire W13247;
wire W13248;
wire W13249;
wire W13250;
wire W13251;
wire W13252;
wire W13253;
wire W13254;
wire W13255;
wire W13256;
wire W13257;
wire W13258;
wire W13259;
wire W13260;
wire W13261;
wire W13262;
wire W13263;
wire W13264;
wire W13265;
wire W13266;
wire W13267;
wire W13268;
wire W13269;
wire W13270;
wire W13271;
wire W13272;
wire W13273;
wire W13274;
wire W13275;
wire W13276;
wire W13277;
wire W13278;
wire W13279;
wire W13280;
wire W13281;
wire W13282;
wire W13283;
wire W13284;
wire W13285;
wire W13286;
wire W13287;
wire W13288;
wire W13289;
wire W13290;
wire W13291;
wire W13292;
wire W13293;
wire W13294;
wire W13295;
wire W13296;
wire W13297;
wire W13298;
wire W13299;
wire W13300;
wire W13301;
wire W13302;
wire W13303;
wire W13304;
wire W13305;
wire W13306;
wire W13307;
wire W13308;
wire W13309;
wire W13310;
wire W13311;
wire W13312;
wire W13313;
wire W13314;
wire W13315;
wire W13316;
wire W13317;
wire W13318;
wire W13319;
wire W13320;
wire W13321;
wire W13322;
wire W13323;
wire W13324;
wire W13325;
wire W13326;
wire W13327;
wire W13328;
wire W13329;
wire W13330;
wire W13331;
wire W13332;
wire W13333;
wire W13334;
wire W13335;
wire W13336;
wire W13337;
wire W13338;
wire W13339;
wire W13340;
wire W13341;
wire W13342;
wire W13343;
wire W13344;
wire W13345;
wire W13346;
wire W13347;
wire W13348;
wire W13349;
wire W13350;
wire W13351;
wire W13352;
wire W13353;
wire W13354;
wire W13355;
wire W13356;
wire W13357;
wire W13358;
wire W13359;
wire W13360;
wire W13361;
wire W13362;
wire W13363;
wire W13364;
wire W13365;
wire W13366;
wire W13367;
wire W13368;
wire W13369;
wire W13370;
wire W13371;
wire W13372;
wire W13373;
wire W13374;
wire W13375;
wire W13376;
wire W13377;
wire W13378;
wire W13379;
wire W13380;
wire W13381;
wire W13382;
wire W13383;
wire W13384;
wire W13385;
wire W13386;
wire W13387;
wire W13388;
wire W13389;
wire W13390;
wire W13391;
wire W13392;
wire W13393;
wire W13394;
wire W13395;
wire W13396;
wire W13397;
wire W13398;
wire W13399;
wire W13400;
wire W13401;
wire W13402;
wire W13403;
wire W13404;
wire W13405;
wire W13406;
wire W13407;
wire W13408;
wire W13409;
wire W13410;
wire W13411;
wire W13412;
wire W13413;
wire W13414;
wire W13415;
wire W13416;
wire W13417;
wire W13418;
wire W13419;
wire W13420;
wire W13421;
wire W13422;
wire W13423;
wire W13424;
wire W13425;
wire W13426;
wire W13427;
wire W13428;
wire W13429;
wire W13430;
wire W13431;
wire W13432;
wire W13433;
wire W13434;
wire W13435;
wire W13436;
wire W13437;
wire W13438;
wire W13439;
wire W13440;
wire W13441;
wire W13442;
wire W13443;
wire W13444;
wire W13445;
wire W13446;
wire W13447;
wire W13448;
wire W13449;
wire W13450;
wire W13451;
wire W13452;
wire W13453;
wire W13454;
wire W13455;
wire W13456;
wire W13457;
wire W13458;
wire W13459;
wire W13460;
wire W13461;
wire W13462;
wire W13463;
wire W13464;
wire W13465;
wire W13466;
wire W13467;
wire W13468;
wire W13469;
wire W13470;
wire W13471;
wire W13472;
wire W13473;
wire W13474;
wire W13475;
wire W13476;
wire W13477;
wire W13478;
wire W13479;
wire W13480;
wire W13481;
wire W13482;
wire W13483;
wire W13484;
wire W13485;
wire W13486;
wire W13487;
wire W13488;
wire W13489;
wire W13490;
wire W13491;
wire W13492;
wire W13493;
wire W13494;
wire W13495;
wire W13496;
wire W13497;
wire W13498;
wire W13499;
wire W13500;
wire W13501;
wire W13502;
wire W13503;
wire W13504;
wire W13505;
wire W13506;
wire W13507;
wire W13508;
wire W13509;
wire W13510;
wire W13511;
wire W13512;
wire W13513;
wire W13514;
wire W13515;
wire W13516;
wire W13517;
wire W13518;
wire W13519;
wire W13520;
wire W13521;
wire W13522;
wire W13523;
wire W13524;
wire W13525;
wire W13526;
wire W13527;
wire W13528;
wire W13529;
wire W13530;
wire W13531;
wire W13532;
wire W13533;
wire W13534;
wire W13535;
wire W13536;
wire W13537;
wire W13538;
wire W13539;
wire W13540;
wire W13541;
wire W13542;
wire W13543;
wire W13544;
wire W13545;
wire W13546;
wire W13547;
wire W13548;
wire W13549;
wire W13550;
wire W13551;
wire W13552;
wire W13553;
wire W13554;
wire W13555;
wire W13556;
wire W13557;
wire W13558;
wire W13559;
wire W13560;
wire W13561;
wire W13562;
wire W13563;
wire W13564;
wire W13565;
wire W13566;
wire W13567;
wire W13568;
wire W13569;
wire W13570;
wire W13571;
wire W13572;
wire W13573;
wire W13574;
wire W13575;
wire W13576;
wire W13577;
wire W13578;
wire W13579;
wire W13580;
wire W13581;
wire W13582;
wire W13583;
wire W13584;
wire W13585;
wire W13586;
wire W13587;
wire W13588;
wire W13589;
wire W13590;
wire W13591;
wire W13592;
wire W13593;
wire W13594;
wire W13595;
wire W13596;
wire W13597;
wire W13598;
wire W13599;
wire W13600;
wire W13601;
wire W13602;
wire W13603;
wire W13604;
wire W13605;
wire W13606;
wire W13607;
wire W13608;
wire W13609;
wire W13610;
wire W13611;
wire W13612;
wire W13613;
wire W13614;
wire W13615;
wire W13616;
wire W13617;
wire W13618;
wire W13619;
wire W13620;
wire W13621;
wire W13622;
wire W13623;
wire W13624;
wire W13625;
wire W13626;
wire W13627;
wire W13628;
wire W13629;
wire W13630;
wire W13631;
wire W13632;
wire W13633;
wire W13634;
wire W13635;
wire W13636;
wire W13637;
wire W13638;
wire W13639;
wire W13640;
wire W13641;
wire W13642;
wire W13643;
wire W13644;
wire W13645;
wire W13646;
wire W13647;
wire W13648;
wire W13649;
wire W13650;
wire W13651;
wire W13652;
wire W13653;
wire W13654;
wire W13655;
wire W13656;
wire W13657;
wire W13658;
wire W13659;
wire W13660;
wire W13661;
wire W13662;
wire W13663;
wire W13664;
wire W13665;
wire W13666;
wire W13667;
wire W13668;
wire W13669;
wire W13670;
wire W13671;
wire W13672;
wire W13673;
wire W13674;
wire W13675;
wire W13676;
wire W13677;
wire W13678;
wire W13679;
wire W13680;
wire W13681;
wire W13682;
wire W13683;
wire W13684;
wire W13685;
wire W13686;
wire W13687;
wire W13688;
wire W13689;
wire W13690;
wire W13691;
wire W13692;
wire W13693;
wire W13694;
wire W13695;
wire W13696;
wire W13697;
wire W13698;
wire W13699;
wire W13700;
wire W13701;
wire W13702;
wire W13703;
wire W13704;
wire W13705;
wire W13706;
wire W13707;
wire W13708;
wire W13709;
wire W13710;
wire W13711;
wire W13712;
wire W13713;
wire W13714;
wire W13715;
wire W13716;
wire W13717;
wire W13718;
wire W13719;
wire W13720;
wire W13721;
wire W13722;
wire W13723;
wire W13724;
wire W13725;
wire W13726;
wire W13727;
wire W13728;
wire W13729;
wire W13730;
wire W13731;
wire W13732;
wire W13733;
wire W13734;
wire W13735;
wire W13736;
wire W13737;
wire W13738;
wire W13739;
wire W13740;
wire W13741;
wire W13742;
wire W13743;
wire W13744;
wire W13745;
wire W13746;
wire W13747;
wire W13748;
wire W13749;
wire W13750;
wire W13751;
wire W13752;
wire W13753;
wire W13754;
wire W13755;
wire W13756;
wire W13757;
wire W13758;
wire W13759;
wire W13760;
wire W13761;
wire W13762;
wire W13763;
wire W13764;
wire W13765;
wire W13766;
wire W13767;
wire W13768;
wire W13769;
wire W13770;
wire W13771;
wire W13772;
wire W13773;
wire W13774;
wire W13775;
wire W13776;
wire W13777;
wire W13778;
wire W13779;
wire W13780;
wire W13781;
wire W13782;
wire W13783;
wire W13784;
wire W13785;
wire W13786;
wire W13787;
wire W13788;
wire W13789;
wire W13790;
wire W13791;
wire W13792;
wire W13793;
wire W13794;
wire W13795;
wire W13796;
wire W13797;
wire W13798;
wire W13799;
wire W13800;
wire W13801;
wire W13802;
wire W13803;
wire W13804;
wire W13805;
wire W13806;
wire W13807;
wire W13808;
wire W13809;
wire W13810;
wire W13811;
wire W13812;
wire W13813;
wire W13814;
wire W13815;
wire W13816;
wire W13817;
wire W13818;
wire W13819;
wire W13820;
wire W13821;
wire W13822;
wire W13823;
wire W13824;
wire W13825;
wire W13826;
wire W13827;
wire W13828;
wire W13829;
wire W13830;
wire W13831;
wire W13832;
wire W13833;
wire W13834;
wire W13835;
wire W13836;
wire W13837;
wire W13838;
wire W13839;
wire W13840;
wire W13841;
wire W13842;
wire W13843;
wire W13844;
wire W13845;
wire W13846;
wire W13847;
wire W13848;
wire W13849;
wire W13850;
wire W13851;
wire W13852;
wire W13853;
wire W13854;
wire W13855;
wire W13856;
wire W13857;
wire W13858;
wire W13859;
wire W13860;
wire W13861;
wire W13862;
wire W13863;
wire W13864;
wire W13865;
wire W13866;
wire W13867;
wire W13868;
wire W13869;
wire W13870;
wire W13871;
wire W13872;
wire W13873;
wire W13874;
wire W13875;
wire W13876;
wire W13877;
wire W13878;
wire W13879;
wire W13880;
wire W13881;
wire W13882;
wire W13883;
wire W13884;
wire W13885;
wire W13886;
wire W13887;
wire W13888;
wire W13889;
wire W13890;
wire W13891;
wire W13892;
wire W13893;
wire W13894;
wire W13895;
wire W13896;
wire W13897;
wire W13898;
wire W13899;
wire W13900;
wire W13901;
wire W13902;
wire W13903;
wire W13904;
wire W13905;
wire W13906;
wire W13907;
wire W13908;
wire W13909;
wire W13910;
wire W13911;
wire W13912;
wire W13913;
wire W13914;
wire W13915;
wire W13916;
wire W13917;
wire W13918;
wire W13919;
wire W13920;
wire W13921;
wire W13922;
wire W13923;
wire W13924;
wire W13925;
wire W13926;
wire W13927;
wire W13928;
wire W13929;
wire W13930;
wire W13931;
wire W13932;
wire W13933;
wire W13934;
wire W13935;
wire W13936;
wire W13937;
wire W13938;
wire W13939;
wire W13940;
wire W13941;
wire W13942;
wire W13943;
wire W13944;
wire W13945;
wire W13946;
wire W13947;
wire W13948;
wire W13949;
wire W13950;
wire W13951;
wire W13952;
wire W13953;
wire W13954;
wire W13955;
wire W13956;
wire W13957;
wire W13958;
wire W13959;
wire W13960;
wire W13961;
wire W13962;
wire W13963;
wire W13964;
wire W13965;
wire W13966;
wire W13967;
wire W13968;
wire W13969;
wire W13970;
wire W13971;
wire W13972;
wire W13973;
wire W13974;
wire W13975;
wire W13976;
wire W13977;
wire W13978;
wire W13979;
wire W13980;
wire W13981;
wire W13982;
wire W13983;
wire W13984;
wire W13985;
wire W13986;
wire W13987;
wire W13988;
wire W13989;
wire W13990;
wire W13991;
wire W13992;
wire W13993;
wire W13994;
wire W13995;
wire W13996;
wire W13997;
wire W13998;
wire W13999;
wire W14000;
wire W14001;
wire W14002;
wire W14003;
wire W14004;
wire W14005;
wire W14006;
wire W14007;
wire W14008;
wire W14009;
wire W14010;
wire W14011;
wire W14012;
wire W14013;
wire W14014;
wire W14015;
wire W14016;
wire W14017;
wire W14018;
wire W14019;
wire W14020;
wire W14021;
wire W14022;
wire W14023;
wire W14024;
wire W14025;
wire W14026;
wire W14027;
wire W14028;
wire W14029;
wire W14030;
wire W14031;
wire W14032;
wire W14033;
wire W14034;
wire W14035;
wire W14036;
wire W14037;
wire W14038;
wire W14039;
wire W14040;
wire W14041;
wire W14042;
wire W14043;
wire W14044;
wire W14045;
wire W14046;
wire W14047;
wire W14048;
wire W14049;
wire W14050;
wire W14051;
wire W14052;
wire W14053;
wire W14054;
wire W14055;
wire W14056;
wire W14057;
wire W14058;
wire W14059;
wire W14060;
wire W14061;
wire W14062;
wire W14063;
wire W14064;
wire W14065;
wire W14066;
wire W14067;
wire W14068;
wire W14069;
wire W14070;
wire W14071;
wire W14072;
wire W14073;
wire W14074;
wire W14075;
wire W14076;
wire W14077;
wire W14078;
wire W14079;
wire W14080;
wire W14081;
wire W14082;
wire W14083;
wire W14084;
wire W14085;
wire W14086;
wire W14087;
wire W14088;
wire W14089;
wire W14090;
wire W14091;
wire W14092;
wire W14093;
wire W14094;
wire W14095;
wire W14096;
wire W14097;
wire W14098;
wire W14099;
wire W14100;
wire W14101;
wire W14102;
wire W14103;
wire W14104;
wire W14105;
wire W14106;
wire W14107;
wire W14108;
wire W14109;
wire W14110;
wire W14111;
wire W14112;
wire W14113;
wire W14114;
wire W14115;
wire W14116;
wire W14117;
wire W14118;
wire W14119;
wire W14120;
wire W14121;
wire W14122;
wire W14123;
wire W14124;
wire W14125;
wire W14126;
wire W14127;
wire W14128;
wire W14129;
wire W14130;
wire W14131;
wire W14132;
wire W14133;
wire W14134;
wire W14135;
wire W14136;
wire W14137;
wire W14138;
wire W14139;
wire W14140;
wire W14141;
wire W14142;
wire W14143;
wire W14144;
wire W14145;
wire W14146;
wire W14147;
wire W14148;
wire W14149;
wire W14150;
wire W14151;
wire W14152;
wire W14153;
wire W14154;
wire W14155;
wire W14156;
wire W14157;
wire W14158;
wire W14159;
wire W14160;
wire W14161;
wire W14162;
wire W14163;
wire W14164;
wire W14165;
wire W14166;
wire W14167;
wire W14168;
wire W14169;
wire W14170;
wire W14171;
wire W14172;
wire W14173;
wire W14174;
wire W14175;
wire W14176;
wire W14177;
wire W14178;
wire W14179;
wire W14180;
wire W14181;
wire W14182;
wire W14183;
wire W14184;
wire W14185;
wire W14186;
wire W14187;
wire W14188;
wire W14189;
wire W14190;
wire W14191;
wire W14192;
wire W14193;
wire W14194;
wire W14195;
wire W14196;
wire W14197;
wire W14198;
wire W14199;
wire W14200;
wire W14201;
wire W14202;
wire W14203;
wire W14204;
wire W14205;
wire W14206;
wire W14207;
wire W14208;
wire W14209;
wire W14210;
wire W14211;
wire W14212;
wire W14213;
wire W14214;
wire W14215;
wire W14216;
wire W14217;
wire W14218;
wire W14219;
wire W14220;
wire W14221;
wire W14222;
wire W14223;
wire W14224;
wire W14225;
wire W14226;
wire W14227;
wire W14228;
wire W14229;
wire W14230;
wire W14231;
wire W14232;
wire W14233;
wire W14234;
wire W14235;
wire W14236;
wire W14237;
wire W14238;
wire W14239;
wire W14240;
wire W14241;
wire W14242;
wire W14243;
wire W14244;
wire W14245;
wire W14246;
wire W14247;
wire W14248;
wire W14249;
wire W14250;
wire W14251;
wire W14252;
wire W14253;
wire W14254;
wire W14255;
wire W14256;
wire W14257;
wire W14258;
wire W14259;
wire W14260;
wire W14261;
wire W14262;
wire W14263;
wire W14264;
wire W14265;
wire W14266;
wire W14267;
wire W14268;
wire W14269;
wire W14270;
wire W14271;
wire W14272;
wire W14273;
wire W14274;
wire W14275;
wire W14276;
wire W14277;
wire W14278;
wire W14279;
wire W14280;
wire W14281;
wire W14282;
wire W14283;
wire W14284;
wire W14285;
wire W14286;
wire W14287;
wire W14288;
wire W14289;
wire W14290;
wire W14291;
wire W14292;
wire W14293;
wire W14294;
wire W14295;
wire W14296;
wire W14297;
wire W14298;
wire W14299;
wire W14300;
wire W14301;
wire W14302;
wire W14303;
wire W14304;
wire W14305;
wire W14306;
wire W14307;
wire W14308;
wire W14309;
wire W14310;
wire W14311;
wire W14312;
wire W14313;
wire W14314;
wire W14315;
wire W14316;
wire W14317;
wire W14318;
wire W14319;
wire W14320;
wire W14321;
wire W14322;
wire W14323;
wire W14324;
wire W14325;
wire W14326;
wire W14327;
wire W14328;
wire W14329;
wire W14330;
wire W14331;
wire W14332;
wire W14333;
wire W14334;
wire W14335;
wire W14336;
wire W14337;
wire W14338;
wire W14339;
wire W14340;
wire W14341;
wire W14342;
wire W14343;
wire W14344;
wire W14345;
wire W14346;
wire W14347;
wire W14348;
wire W14349;
wire W14350;
wire W14351;
wire W14352;
wire W14353;
wire W14354;
wire W14355;
wire W14356;
wire W14357;
wire W14358;
wire W14359;
wire W14360;
wire W14361;
wire W14362;
wire W14363;
wire W14364;
wire W14365;
wire W14366;
wire W14367;
wire W14368;
wire W14369;
wire W14370;
wire W14371;
wire W14372;
wire W14373;
wire W14374;
wire W14375;
wire W14376;
wire W14377;
wire W14378;
wire W14379;
wire W14380;
wire W14381;
wire W14382;
wire W14383;
wire W14384;
wire W14385;
wire W14386;
wire W14387;
wire W14388;
wire W14389;
wire W14390;
wire W14391;
wire W14392;
wire W14393;
wire W14394;
wire W14395;
wire W14396;
wire W14397;
wire W14398;
wire W14399;
wire W14400;
wire W14401;
wire W14402;
wire W14403;
wire W14404;
wire W14405;
wire W14406;
wire W14407;
wire W14408;
wire W14409;
wire W14410;
wire W14411;
wire W14412;
wire W14413;
wire W14414;
wire W14415;
wire W14416;
wire W14417;
wire W14418;
wire W14419;
wire W14420;
wire W14421;
wire W14422;
wire W14423;
wire W14424;
wire W14425;
wire W14426;
wire W14427;
wire W14428;
wire W14429;
wire W14430;
wire W14431;
wire W14432;
wire W14433;
wire W14434;
wire W14435;
wire W14436;
wire W14437;
wire W14438;
wire W14439;
wire W14440;
wire W14441;
wire W14442;
wire W14443;
wire W14444;
wire W14445;
wire W14446;
wire W14447;
wire W14448;
wire W14449;
wire W14450;
wire W14451;
wire W14452;
wire W14453;
wire W14454;
wire W14455;
wire W14456;
wire W14457;
wire W14458;
wire W14459;
wire W14460;
wire W14461;
wire W14462;
wire W14463;
wire W14464;
wire W14465;
wire W14466;
wire W14467;
wire W14468;
wire W14469;
wire W14470;
wire W14471;
wire W14472;
wire W14473;
wire W14474;
wire W14475;
wire W14476;
wire W14477;
wire W14478;
wire W14479;
wire W14480;
wire W14481;
wire W14482;
wire W14483;
wire W14484;
wire W14485;
wire W14486;
wire W14487;
wire W14488;
wire W14489;
wire W14490;
wire W14491;
wire W14492;
wire W14493;
wire W14494;
wire W14495;
wire W14496;
wire W14497;
wire W14498;
wire W14499;
wire W14500;
wire W14501;
wire W14502;
wire W14503;
wire W14504;
wire W14505;
wire W14506;
wire W14507;
wire W14508;
wire W14509;
wire W14510;
wire W14511;
wire W14512;
wire W14513;
wire W14514;
wire W14515;
wire W14516;
wire W14517;
wire W14518;
wire W14519;
wire W14520;
wire W14521;
wire W14522;
wire W14523;
wire W14524;
wire W14525;
wire W14526;
wire W14527;
wire W14528;
wire W14529;
wire W14530;
wire W14531;
wire W14532;
wire W14533;
wire W14534;
wire W14535;
wire W14536;
wire W14537;
wire W14538;
wire W14539;
wire W14540;
wire W14541;
wire W14542;
wire W14543;
wire W14544;
wire W14545;
wire W14546;
wire W14547;
wire W14548;
wire W14549;
wire W14550;
wire W14551;
wire W14552;
wire W14553;
wire W14554;
wire W14555;
wire W14556;
wire W14557;
wire W14558;
wire W14559;
wire W14560;
wire W14561;
wire W14562;
wire W14563;
wire W14564;
wire W14565;
wire W14566;
wire W14567;
wire W14568;
wire W14569;
wire W14570;
wire W14571;
wire W14572;
wire W14573;
wire W14574;
wire W14575;
wire W14576;
wire W14577;
wire W14578;
wire W14579;
wire W14580;
wire W14581;
wire W14582;
wire W14583;
wire W14584;
wire W14585;
wire W14586;
wire W14587;
wire W14588;
wire W14589;
wire W14590;
wire W14591;
wire W14592;
wire W14593;
wire W14594;
wire W14595;
wire W14596;
wire W14597;
wire W14598;
wire W14599;
wire W14600;
wire W14601;
wire W14602;
wire W14603;
wire W14604;
wire W14605;
wire W14606;
wire W14607;
wire W14608;
wire W14609;
wire W14610;
wire W14611;
wire W14612;
wire W14613;
wire W14614;
wire W14615;
wire W14616;
wire W14617;
wire W14618;
wire W14619;
wire W14620;
wire W14621;
wire W14622;
wire W14623;
wire W14624;
wire W14625;
wire W14626;
wire W14627;
wire W14628;
wire W14629;
wire W14630;
wire W14631;
wire W14632;
wire W14633;
wire W14634;
wire W14635;
wire W14636;
wire W14637;
wire W14638;
wire W14639;
wire W14640;
wire W14641;
wire W14642;
wire W14643;
wire W14644;
wire W14645;
wire W14646;
wire W14647;
wire W14648;
wire W14649;
wire W14650;
wire W14651;
wire W14652;
wire W14653;
wire W14654;
wire W14655;
wire W14656;
wire W14657;
wire W14658;
wire W14659;
wire W14660;
wire W14661;
wire W14662;
wire W14663;
wire W14664;
wire W14665;
wire W14666;
wire W14667;
wire W14668;
wire W14669;
wire W14670;
wire W14671;
wire W14672;
wire W14673;
wire W14674;
wire W14675;
wire W14676;
wire W14677;
wire W14678;
wire W14679;
wire W14680;
wire W14681;
wire W14682;
wire W14683;
wire W14684;
wire W14685;
wire W14686;
wire W14687;
wire W14688;
wire W14689;
wire W14690;
wire W14691;
wire W14692;
wire W14693;
wire W14694;
wire W14695;
wire W14696;
wire W14697;
wire W14698;
wire W14699;
wire W14700;
wire W14701;
wire W14702;
wire W14703;
wire W14704;
wire W14705;
wire W14706;
wire W14707;
wire W14708;
wire W14709;
wire W14710;
wire W14711;
wire W14712;
wire W14713;
wire W14714;
wire W14715;
wire W14716;
wire W14717;
wire W14718;
wire W14719;
wire W14720;
wire W14721;
wire W14722;
wire W14723;
wire W14724;
wire W14725;
wire W14726;
wire W14727;
wire W14728;
wire W14729;
wire W14730;
wire W14731;
wire W14732;
wire W14733;
wire W14734;
wire W14735;
wire W14736;
wire W14737;
wire W14738;
wire W14739;
wire W14740;
wire W14741;
wire W14742;
wire W14743;
wire W14744;
wire W14745;
wire W14746;
wire W14747;
wire W14748;
wire W14749;
wire W14750;
wire W14751;
wire W14752;
wire W14753;
wire W14754;
wire W14755;
wire W14756;
wire W14757;
wire W14758;
wire W14759;
wire W14760;
wire W14761;
wire W14762;
wire W14763;
wire W14764;
wire W14765;
wire W14766;
wire W14767;
wire W14768;
wire W14769;
wire W14770;
wire W14771;
wire W14772;
wire W14773;
wire W14774;
wire W14775;
wire W14776;
wire W14777;
wire W14778;
wire W14779;
wire W14780;
wire W14781;
wire W14782;
wire W14783;
wire W14784;
wire W14785;
wire W14786;
wire W14787;
wire W14788;
wire W14789;
wire W14790;
wire W14791;
wire W14792;
wire W14793;
wire W14794;
wire W14795;
wire W14796;
wire W14797;
wire W14798;
wire W14799;
wire W14800;
wire W14801;
wire W14802;
wire W14803;
wire W14804;
wire W14805;
wire W14806;
wire W14807;
wire W14808;
wire W14809;
wire W14810;
wire W14811;
wire W14812;
wire W14813;
wire W14814;
wire W14815;
wire W14816;
wire W14817;
wire W14818;
wire W14819;
wire W14820;
wire W14821;
wire W14822;
wire W14823;
wire W14824;
wire W14825;
wire W14826;
wire W14827;
wire W14828;
wire W14829;
wire W14830;
wire W14831;
wire W14832;
wire W14833;
wire W14834;
wire W14835;
wire W14836;
wire W14837;
wire W14838;
wire W14839;
wire W14840;
wire W14841;
wire W14842;
wire W14843;
wire W14844;
wire W14845;
wire W14846;
wire W14847;
wire W14848;
wire W14849;
wire W14850;
wire W14851;
wire W14852;
wire W14853;
wire W14854;
wire W14855;
wire W14856;
wire W14857;
wire W14858;
wire W14859;
wire W14860;
wire W14861;
wire W14862;
wire W14863;
wire W14864;
wire W14865;
wire W14866;
wire W14867;
wire W14868;
wire W14869;
wire W14870;
wire W14871;
wire W14872;
wire W14873;
wire W14874;
wire W14875;
wire W14876;
wire W14877;
wire W14878;
wire W14879;
wire W14880;
wire W14881;
wire W14882;
wire W14883;
wire W14884;
wire W14885;
wire W14886;
wire W14887;
wire W14888;
wire W14889;
wire W14890;
wire W14891;
wire W14892;
wire W14893;
wire W14894;
wire W14895;
wire W14896;
wire W14897;
wire W14898;
wire W14899;
wire W14900;
wire W14901;
wire W14902;
wire W14903;
wire W14904;
wire W14905;
wire W14906;
wire W14907;
wire W14908;
wire W14909;
wire W14910;
wire W14911;
wire W14912;
wire W14913;
wire W14914;
wire W14915;
wire W14916;
wire W14917;
wire W14918;
wire W14919;
wire W14920;
wire W14921;
wire W14922;
wire W14923;
wire W14924;
wire W14925;
wire W14926;
wire W14927;
wire W14928;
wire W14929;
wire W14930;
wire W14931;
wire W14932;
wire W14933;
wire W14934;
wire W14935;
wire W14936;
wire W14937;
wire W14938;
wire W14939;
wire W14940;
wire W14941;
wire W14942;
wire W14943;
wire W14944;
wire W14945;
wire W14946;
wire W14947;
wire W14948;
wire W14949;
wire W14950;
wire W14951;
wire W14952;
wire W14953;
wire W14954;
wire W14955;
wire W14956;
wire W14957;
wire W14958;
wire W14959;
wire W14960;
wire W14961;
wire W14962;
wire W14963;
wire W14964;
wire W14965;
wire W14966;
wire W14967;
wire W14968;
wire W14969;
wire W14970;
wire W14971;
wire W14972;
wire W14973;
wire W14974;
wire W14975;
wire W14976;
wire W14977;
wire W14978;
wire W14979;
wire W14980;
wire W14981;
wire W14982;
wire W14983;
wire W14984;
wire W14985;
wire W14986;
wire W14987;
wire W14988;
wire W14989;
wire W14990;
wire W14991;
wire W14992;
wire W14993;
wire W14994;
wire W14995;
wire W14996;
wire W14997;
wire W14998;
wire W14999;
wire W15000;
wire W15001;
wire W15002;
wire W15003;
wire W15004;
wire W15005;
wire W15006;
wire W15007;
wire W15008;
wire W15009;
wire W15010;
wire W15011;
wire W15012;
wire W15013;
wire W15014;
wire W15015;
wire W15016;
wire W15017;
wire W15018;
wire W15019;
wire W15020;
wire W15021;
wire W15022;
wire W15023;
wire W15024;
wire W15025;
wire W15026;
wire W15027;
wire W15028;
wire W15029;
wire W15030;
wire W15031;
wire W15032;
wire W15033;
wire W15034;
wire W15035;
wire W15036;
wire W15037;
wire W15038;
wire W15039;
wire W15040;
wire W15041;
wire W15042;
wire W15043;
wire W15044;
wire W15045;
wire W15046;
wire W15047;
wire W15048;
wire W15049;
wire W15050;
wire W15051;
wire W15052;
wire W15053;
wire W15054;
wire W15055;
wire W15056;
wire W15057;
wire W15058;
wire W15059;
wire W15060;
wire W15061;
wire W15062;
wire W15063;
wire W15064;
wire W15065;
wire W15066;
wire W15067;
wire W15068;
wire W15069;
wire W15070;
wire W15071;
wire W15072;
wire W15073;
wire W15074;
wire W15075;
wire W15076;
wire W15077;
wire W15078;
wire W15079;
wire W15080;
wire W15081;
wire W15082;
wire W15083;
wire W15084;
wire W15085;
wire W15086;
wire W15087;
wire W15088;
wire W15089;
wire W15090;
wire W15091;
wire W15092;
wire W15093;
wire W15094;
wire W15095;
wire W15096;
wire W15097;
wire W15098;
wire W15099;
wire W15100;
wire W15101;
wire W15102;
wire W15103;
wire W15104;
wire W15105;
wire W15106;
wire W15107;
wire W15108;
wire W15109;
wire W15110;
wire W15111;
wire W15112;
wire W15113;
wire W15114;
wire W15115;
wire W15116;
wire W15117;
wire W15118;
wire W15119;
wire W15120;
wire W15121;
wire W15122;
wire W15123;
wire W15124;
wire W15125;
wire W15126;
wire W15127;
wire W15128;
wire W15129;
wire W15130;
wire W15131;
wire W15132;
wire W15133;
wire W15134;
wire W15135;
wire W15136;
wire W15137;
wire W15138;
wire W15139;
wire W15140;
wire W15141;
wire W15142;
wire W15143;
wire W15144;
wire W15145;
wire W15146;
wire W15147;
wire W15148;
wire W15149;
wire W15150;
wire W15151;
wire W15152;
wire W15153;
wire W15154;
wire W15155;
wire W15156;
wire W15157;
wire W15158;
wire W15159;
wire W15160;
wire W15161;
wire W15162;
wire W15163;
wire W15164;
wire W15165;
wire W15166;
wire W15167;
wire W15168;
wire W15169;
wire W15170;
wire W15171;
wire W15172;
wire W15173;
wire W15174;
wire W15175;
wire W15176;
wire W15177;
wire W15178;
wire W15179;
wire W15180;
wire W15181;
wire W15182;
wire W15183;
wire W15184;
wire W15185;
wire W15186;
wire W15187;
wire W15188;
wire W15189;
wire W15190;
wire W15191;
wire W15192;
wire W15193;
wire W15194;
wire W15195;
wire W15196;
wire W15197;
wire W15198;
wire W15199;
wire W15200;
wire W15201;
wire W15202;
wire W15203;
wire W15204;
wire W15205;
wire W15206;
wire W15207;
wire W15208;
wire W15209;
wire W15210;
wire W15211;
wire W15212;
wire W15213;
wire W15214;
wire W15215;
wire W15216;
wire W15217;
wire W15218;
wire W15219;
wire W15220;
wire W15221;
wire W15222;
wire W15223;
wire W15224;
wire W15225;
wire W15226;
wire W15227;
wire W15228;
wire W15229;
wire W15230;
wire W15231;
wire W15232;
wire W15233;
wire W15234;
wire W15235;
wire W15236;
wire W15237;
wire W15238;
wire W15239;
wire W15240;
wire W15241;
wire W15242;
wire W15243;
wire W15244;
wire W15245;
wire W15246;
wire W15247;
wire W15248;
wire W15249;
wire W15250;
wire W15251;
wire W15252;
wire W15253;
wire W15254;
wire W15255;
wire W15256;
wire W15257;
wire W15258;
wire W15259;
wire W15260;
wire W15261;
wire W15262;
wire W15263;
wire W15264;
wire W15265;
wire W15266;
wire W15267;
wire W15268;
wire W15269;
wire W15270;
wire W15271;
wire W15272;
wire W15273;
wire W15274;
wire W15275;
wire W15276;
wire W15277;
wire W15278;
wire W15279;
wire W15280;
wire W15281;
wire W15282;
wire W15283;
wire W15284;
wire W15285;
wire W15286;
wire W15287;
wire W15288;
wire W15289;
wire W15290;
wire W15291;
wire W15292;
wire W15293;
wire W15294;
wire W15295;
wire W15296;
wire W15297;
wire W15298;
wire W15299;
wire W15300;
wire W15301;
wire W15302;
wire W15303;
wire W15304;
wire W15305;
wire W15306;
wire W15307;
wire W15308;
wire W15309;
wire W15310;
wire W15311;
wire W15312;
wire W15313;
wire W15314;
wire W15315;
wire W15316;
wire W15317;
wire W15318;
wire W15319;
wire W15320;
wire W15321;
wire W15322;
wire W15323;
wire W15324;
wire W15325;
wire W15326;
wire W15327;
wire W15328;
wire W15329;
wire W15330;
wire W15331;
wire W15332;
wire W15333;
wire W15334;
wire W15335;
wire W15336;
wire W15337;
wire W15338;
wire W15339;
wire W15340;
wire W15341;
wire W15342;
wire W15343;
wire W15344;
wire W15345;
wire W15346;
wire W15347;
wire W15348;
wire W15349;
wire W15350;
wire W15351;
wire W15352;
wire W15353;
wire W15354;
wire W15355;
wire W15356;
wire W15357;
wire W15358;
wire W15359;
wire W15360;
wire W15361;
wire W15362;
wire W15363;
wire W15364;
wire W15365;
wire W15366;
wire W15367;
wire W15368;
wire W15369;
wire W15370;
wire W15371;
wire W15372;
wire W15373;
wire W15374;
wire W15375;
wire W15376;
wire W15377;
wire W15378;
wire W15379;
wire W15380;
wire W15381;
wire W15382;
wire W15383;
wire W15384;
wire W15385;
wire W15386;
wire W15387;
wire W15388;
wire W15389;
wire W15390;
wire W15391;
wire W15392;
wire W15393;
wire W15394;
wire W15395;
wire W15396;
wire W15397;
wire W15398;
wire W15399;
wire W15400;
wire W15401;
wire W15402;
wire W15403;
wire W15404;
wire W15405;
wire W15406;
wire W15407;
wire W15408;
wire W15409;
wire W15410;
wire W15411;
wire W15412;
wire W15413;
wire W15414;
wire W15415;
wire W15416;
wire W15417;
wire W15418;
wire W15419;
wire W15420;
wire W15421;
wire W15422;
wire W15423;
wire W15424;
wire W15425;
wire W15426;
wire W15427;
wire W15428;
wire W15429;
wire W15430;
wire W15431;
wire W15432;
wire W15433;
wire W15434;
wire W15435;
wire W15436;
wire W15437;
wire W15438;
wire W15439;
wire W15440;
wire W15441;
wire W15442;
wire W15443;
wire W15444;
wire W15445;
wire W15446;
wire W15447;
wire W15448;
wire W15449;
wire W15450;
wire W15451;
wire W15452;
wire W15453;
wire W15454;
wire W15455;
wire W15456;
wire W15457;
wire W15458;
wire W15459;
wire W15460;
wire W15461;
wire W15462;
wire W15463;
wire W15464;
wire W15465;
wire W15466;
wire W15467;
wire W15468;
wire W15469;
wire W15470;
wire W15471;
wire W15472;
wire W15473;
wire W15474;
wire W15475;
wire W15476;
wire W15477;
wire W15478;
wire W15479;
wire W15480;
wire W15481;
wire W15482;
wire W15483;
wire W15484;
wire W15485;
wire W15486;
wire W15487;
wire W15488;
wire W15489;
wire W15490;
wire W15491;
wire W15492;
wire W15493;
wire W15494;
wire W15495;
wire W15496;
wire W15497;
wire W15498;
wire W15499;
wire W15500;
wire W15501;
wire W15502;
wire W15503;
wire W15504;
wire W15505;
wire W15506;
wire W15507;
wire W15508;
wire W15509;
wire W15510;
wire W15511;
wire W15512;
wire W15513;
wire W15514;
wire W15515;
wire W15516;
wire W15517;
wire W15518;
wire W15519;
wire W15520;
wire W15521;
wire W15522;
wire W15523;
wire W15524;
wire W15525;
wire W15526;
wire W15527;
wire W15528;
wire W15529;
wire W15530;
wire W15531;
wire W15532;
wire W15533;
wire W15534;
wire W15535;
wire W15536;
wire W15537;
wire W15538;
wire W15539;
wire W15540;
wire W15541;
wire W15542;
wire W15543;
wire W15544;
wire W15545;
wire W15546;
wire W15547;
wire W15548;
wire W15549;
wire W15550;
wire W15551;
wire W15552;
wire W15553;
wire W15554;
wire W15555;
wire W15556;
wire W15557;
wire W15558;
wire W15559;
wire W15560;
wire W15561;
wire W15562;
wire W15563;
wire W15564;
wire W15565;
wire W15566;
wire W15567;
wire W15568;
wire W15569;
wire W15570;
wire W15571;
wire W15572;
wire W15573;
wire W15574;
wire W15575;
wire W15576;
wire W15577;
wire W15578;
wire W15579;
wire W15580;
wire W15581;
wire W15582;
wire W15583;
wire W15584;
wire W15585;
wire W15586;
wire W15587;
wire W15588;
wire W15589;
wire W15590;
wire W15591;
wire W15592;
wire W15593;
wire W15594;
wire W15595;
wire W15596;
wire W15597;
wire W15598;
wire W15599;
wire W15600;
wire W15601;
wire W15602;
wire W15603;
wire W15604;
wire W15605;
wire W15606;
wire W15607;
wire W15608;
wire W15609;
wire W15610;
wire W15611;
wire W15612;
wire W15613;
wire W15614;
wire W15615;
wire W15616;
wire W15617;
wire W15618;
wire W15619;
wire W15620;
wire W15621;
wire W15622;
wire W15623;
wire W15624;
wire W15625;
wire W15626;
wire W15627;
wire W15628;
wire W15629;
wire W15630;
wire W15631;
wire W15632;
wire W15633;
wire W15634;
wire W15635;
wire W15636;
wire W15637;
wire W15638;
wire W15639;
wire W15640;
wire W15641;
wire W15642;
wire W15643;
wire W15644;
wire W15645;
wire W15646;
wire W15647;
wire W15648;
wire W15649;
wire W15650;
wire W15651;
wire W15652;
wire W15653;
wire W15654;
wire W15655;
wire W15656;
wire W15657;
wire W15658;
wire W15659;
wire W15660;
wire W15661;
wire W15662;
wire W15663;
wire W15664;
wire W15665;
wire W15666;
wire W15667;
wire W15668;
wire W15669;
wire W15670;
wire W15671;
wire W15672;
wire W15673;
wire W15674;
wire W15675;
wire W15676;
wire W15677;
wire W15678;
wire W15679;
wire W15680;
wire W15681;
wire W15682;
wire W15683;
wire W15684;
wire W15685;
wire W15686;
wire W15687;
wire W15688;
wire W15689;
wire W15690;
wire W15691;
wire W15692;
wire W15693;
wire W15694;
wire W15695;
wire W15696;
wire W15697;
wire W15698;
wire W15699;
wire W15700;
wire W15701;
wire W15702;
wire W15703;
wire W15704;
wire W15705;
wire W15706;
wire W15707;
wire W15708;
wire W15709;
wire W15710;
wire W15711;
wire W15712;
wire W15713;
wire W15714;
wire W15715;
wire W15716;
wire W15717;
wire W15718;
wire W15719;
wire W15720;
wire W15721;
wire W15722;
wire W15723;
wire W15724;
wire W15725;
wire W15726;
wire W15727;
wire W15728;
wire W15729;
wire W15730;
wire W15731;
wire W15732;
wire W15733;
wire W15734;
wire W15735;
wire W15736;
wire W15737;
wire W15738;
wire W15739;
wire W15740;
wire W15741;
wire W15742;
wire W15743;
wire W15744;
wire W15745;
wire W15746;
wire W15747;
wire W15748;
wire W15749;
wire W15750;
wire W15751;
wire W15752;
wire W15753;
wire W15754;
wire W15755;
wire W15756;
wire W15757;
wire W15758;
wire W15759;
wire W15760;
wire W15761;
wire W15762;
wire W15763;
wire W15764;
wire W15765;
wire W15766;
wire W15767;
wire W15768;
wire W15769;
wire W15770;
wire W15771;
wire W15772;
wire W15773;
wire W15774;
wire W15775;
wire W15776;
wire W15777;
wire W15778;
wire W15779;
wire W15780;
wire W15781;
wire W15782;
wire W15783;
wire W15784;
wire W15785;
wire W15786;
wire W15787;
wire W15788;
wire W15789;
wire W15790;
wire W15791;
wire W15792;
wire W15793;
wire W15794;
wire W15795;
wire W15796;
wire W15797;
wire W15798;
wire W15799;
wire W15800;
wire W15801;
wire W15802;
wire W15803;
wire W15804;
wire W15805;
wire W15806;
wire W15807;
wire W15808;
wire W15809;
wire W15810;
wire W15811;
wire W15812;
wire W15813;
wire W15814;
wire W15815;
wire W15816;
wire W15817;
wire W15818;
wire W15819;
wire W15820;
wire W15821;
wire W15822;
wire W15823;
wire W15824;
wire W15825;
wire W15826;
wire W15827;
wire W15828;
wire W15829;
wire W15830;
wire W15831;
wire W15832;
wire W15833;
wire W15834;
wire W15835;
wire W15836;
wire W15837;
wire W15838;
wire W15839;
wire W15840;
wire W15841;
wire W15842;
wire W15843;
wire W15844;
wire W15845;
wire W15846;
wire W15847;
wire W15848;
wire W15849;
wire W15850;
wire W15851;
wire W15852;
wire W15853;
wire W15854;
wire W15855;
wire W15856;
wire W15857;
wire W15858;
wire W15859;
wire W15860;
wire W15861;
wire W15862;
wire W15863;
wire W15864;
wire W15865;
wire W15866;
wire W15867;
wire W15868;
wire W15869;
wire W15870;
wire W15871;
wire W15872;
wire W15873;
wire W15874;
wire W15875;
wire W15876;
wire W15877;
wire W15878;
wire W15879;
wire W15880;
wire W15881;
wire W15882;
wire W15883;
wire W15884;
wire W15885;
wire W15886;
wire W15887;
wire W15888;
wire W15889;
wire W15890;
wire W15891;
wire W15892;
wire W15893;
wire W15894;
wire W15895;
wire W15896;
wire W15897;
wire W15898;
wire W15899;
wire W15900;
wire W15901;
wire W15902;
wire W15903;
wire W15904;
wire W15905;
wire W15906;
wire W15907;
wire W15908;
wire W15909;
wire W15910;
wire W15911;
wire W15912;
wire W15913;
wire W15914;
wire W15915;
wire W15916;
wire W15917;
wire W15918;
wire W15919;
wire W15920;
wire W15921;
wire W15922;
wire W15923;
wire W15924;
wire W15925;
wire W15926;
wire W15927;
wire W15928;
wire W15929;
wire W15930;
wire W15931;
wire W15932;
wire W15933;
wire W15934;
wire W15935;
wire W15936;
wire W15937;
wire W15938;
wire W15939;
wire W15940;
wire W15941;
wire W15942;
wire W15943;
wire W15944;
wire W15945;
wire W15946;
wire W15947;
wire W15948;
wire W15949;
wire W15950;
wire W15951;
wire W15952;
wire W15953;
wire W15954;
wire W15955;
wire W15956;
wire W15957;
wire W15958;
wire W15959;
wire W15960;
wire W15961;
wire W15962;
wire W15963;
wire W15964;
wire W15965;
wire W15966;
wire W15967;
wire W15968;
wire W15969;
wire W15970;
wire W15971;
wire W15972;
wire W15973;
wire W15974;
wire W15975;
wire W15976;
wire W15977;
wire W15978;
wire W15979;
wire W15980;
wire W15981;
wire W15982;
wire W15983;
wire W15984;
wire W15985;
wire W15986;
wire W15987;
wire W15988;
wire W15989;
wire W15990;
wire W15991;
wire W15992;
wire W15993;
wire W15994;
wire W15995;
wire W15996;
wire W15997;
wire W15998;
wire W15999;
wire W16000;
wire W16001;
wire W16002;
wire W16003;
wire W16004;
wire W16005;
wire W16006;
wire W16007;
wire W16008;
wire W16009;
wire W16010;
wire W16011;
wire W16012;
wire W16013;
wire W16014;
wire W16015;
wire W16016;
wire W16017;
wire W16018;
wire W16019;
wire W16020;
wire W16021;
wire W16022;
wire W16023;
wire W16024;
wire W16025;
wire W16026;
wire W16027;
wire W16028;
wire W16029;
wire W16030;
wire W16031;
wire W16032;
wire W16033;
wire W16034;
wire W16035;
wire W16036;
wire W16037;
wire W16038;
wire W16039;
wire W16040;
wire W16041;
wire W16042;
wire W16043;
wire W16044;
wire W16045;
wire W16046;
wire W16047;
wire W16048;
wire W16049;
wire W16050;
wire W16051;
wire W16052;
wire W16053;
wire W16054;
wire W16055;
wire W16056;
wire W16057;
wire W16058;
wire W16059;
wire W16060;
wire W16061;
wire W16062;
wire W16063;
wire W16064;
wire W16065;
wire W16066;
wire W16067;
wire W16068;
wire W16069;
wire W16070;
wire W16071;
wire W16072;
wire W16073;
wire W16074;
wire W16075;
wire W16076;
wire W16077;
wire W16078;
wire W16079;
wire W16080;
wire W16081;
wire W16082;
wire W16083;
wire W16084;
wire W16085;
wire W16086;
wire W16087;
wire W16088;
wire W16089;
wire W16090;
wire W16091;
wire W16092;
wire W16093;
wire W16094;
wire W16095;
wire W16096;
wire W16097;
wire W16098;
wire W16099;
wire W16100;
wire W16101;
wire W16102;
wire W16103;
wire W16104;
wire W16105;
wire W16106;
wire W16107;
wire W16108;
wire W16109;
wire W16110;
wire W16111;
wire W16112;
wire W16113;
wire W16114;
wire W16115;
wire W16116;
wire W16117;
wire W16118;
wire W16119;
wire W16120;
wire W16121;
wire W16122;
wire W16123;
wire W16124;
wire W16125;
wire W16126;
wire W16127;
wire W16128;
wire W16129;
wire W16130;
wire W16131;
wire W16132;
wire W16133;
wire W16134;
wire W16135;
wire W16136;
wire W16137;
wire W16138;
wire W16139;
wire W16140;
wire W16141;
wire W16142;
wire W16143;
wire W16144;
wire W16145;
wire W16146;
wire W16147;
wire W16148;
wire W16149;
wire W16150;
wire W16151;
wire W16152;
wire W16153;
wire W16154;
wire W16155;
wire W16156;
wire W16157;
wire W16158;
wire W16159;
wire W16160;
wire W16161;
wire W16162;
wire W16163;
wire W16164;
wire W16165;
wire W16166;
wire W16167;
wire W16168;
wire W16169;
wire W16170;
wire W16171;
wire W16172;
wire W16173;
wire W16174;
wire W16175;
wire W16176;
wire W16177;
wire W16178;
wire W16179;
wire W16180;
wire W16181;
wire W16182;
wire W16183;
wire W16184;
wire W16185;
wire W16186;
wire W16187;
wire W16188;
wire W16189;
wire W16190;
wire W16191;
wire W16192;
wire W16193;
wire W16194;
wire W16195;
wire W16196;
wire W16197;
wire W16198;
wire W16199;
wire W16200;
wire W16201;
wire W16202;
wire W16203;
wire W16204;
wire W16205;
wire W16206;
wire W16207;
wire W16208;
wire W16209;
wire W16210;
wire W16211;
wire W16212;
wire W16213;
wire W16214;
wire W16215;
wire W16216;
wire W16217;
wire W16218;
wire W16219;
wire W16220;
wire W16221;
wire W16222;
wire W16223;
wire W16224;
wire W16225;
wire W16226;
wire W16227;
wire W16228;
wire W16229;
wire W16230;
wire W16231;
wire W16232;
wire W16233;
wire W16234;
wire W16235;
wire W16236;
wire W16237;
wire W16238;
wire W16239;
wire W16240;
wire W16241;
wire W16242;
wire W16243;
wire W16244;
wire W16245;
wire W16246;
wire W16247;
wire W16248;
wire W16249;
wire W16250;
wire W16251;
wire W16252;
wire W16253;
wire W16254;
wire W16255;
wire W16256;
wire W16257;
wire W16258;
wire W16259;
wire W16260;
wire W16261;
wire W16262;
wire W16263;
wire W16264;
wire W16265;
wire W16266;
wire W16267;
wire W16268;
wire W16269;
wire W16270;
wire W16271;
wire W16272;
wire W16273;
wire W16274;
wire W16275;
wire W16276;
wire W16277;
wire W16278;
wire W16279;
wire W16280;
wire W16281;
wire W16282;
wire W16283;
wire W16284;
wire W16285;
wire W16286;
wire W16287;
wire W16288;
wire W16289;
wire W16290;
wire W16291;
wire W16292;
wire W16293;
wire W16294;
wire W16295;
wire W16296;
wire W16297;
wire W16298;
wire W16299;
wire W16300;
wire W16301;
wire W16302;
wire W16303;
wire W16304;
wire W16305;
wire W16306;
wire W16307;
wire W16308;
wire W16309;
wire W16310;
wire W16311;
wire W16312;
wire W16313;
wire W16314;
wire W16315;
wire W16316;
wire W16317;
wire W16318;
wire W16319;
wire W16320;
wire W16321;
wire W16322;
wire W16323;
wire W16324;
wire W16325;
wire W16326;
wire W16327;
wire W16328;
wire W16329;
wire W16330;
wire W16331;
wire W16332;
wire W16333;
wire W16334;
wire W16335;
wire W16336;
wire W16337;
wire W16338;
wire W16339;
wire W16340;
wire W16341;
wire W16342;
wire W16343;
wire W16344;
wire W16345;
wire W16346;
wire W16347;
wire W16348;
wire W16349;
wire W16350;
wire W16351;
wire W16352;
wire W16353;
wire W16354;
wire W16355;
wire W16356;
wire W16357;
wire W16358;
wire W16359;
wire W16360;
wire W16361;
wire W16362;
wire W16363;
wire W16364;
wire W16365;
wire W16366;
wire W16367;
wire W16368;
wire W16369;
wire W16370;
wire W16371;
wire W16372;
wire W16373;
wire W16374;
wire W16375;
wire W16376;
wire W16377;
wire W16378;
wire W16379;
wire W16380;
wire W16381;
wire W16382;
wire W16383;
wire W16384;
wire W16385;
wire W16386;
wire W16387;
wire W16388;
wire W16389;
wire W16390;
wire W16391;
wire W16392;
wire W16393;
wire W16394;
wire W16395;
wire W16396;
wire W16397;
wire W16398;
wire W16399;
wire W16400;
wire W16401;
wire W16402;
wire W16403;
wire W16404;
wire W16405;
wire W16406;
wire W16407;
wire W16408;
wire W16409;
wire W16410;
wire W16411;
wire W16412;
wire W16413;
wire W16414;
wire W16415;
wire W16416;
wire W16417;
wire W16418;
wire W16419;
wire W16420;
wire W16421;
wire W16422;
wire W16423;
wire W16424;
wire W16425;
wire W16426;
wire W16427;
wire W16428;
wire W16429;
wire W16430;
wire W16431;
wire W16432;
wire W16433;
wire W16434;
wire W16435;
wire W16436;
wire W16437;
wire W16438;
wire W16439;
wire W16440;
wire W16441;
wire W16442;
wire W16443;
wire W16444;
wire W16445;
wire W16446;
wire W16447;
wire W16448;
wire W16449;
wire W16450;
wire W16451;
wire W16452;
wire W16453;
wire W16454;
wire W16455;
wire W16456;
wire W16457;
wire W16458;
wire W16459;
wire W16460;
wire W16461;
wire W16462;
wire W16463;
wire W16464;
wire W16465;
wire W16466;
wire W16467;
wire W16468;
wire W16469;
wire W16470;
wire W16471;
wire W16472;
wire W16473;
wire W16474;
wire W16475;
wire W16476;
wire W16477;
wire W16478;
wire W16479;
wire W16480;
wire W16481;
wire W16482;
wire W16483;
wire W16484;
wire W16485;
wire W16486;
wire W16487;
wire W16488;
wire W16489;
wire W16490;
wire W16491;
wire W16492;
wire W16493;
wire W16494;
wire W16495;
wire W16496;
wire W16497;
wire W16498;
wire W16499;
wire W16500;
wire W16501;
wire W16502;
wire W16503;
wire W16504;
wire W16505;
wire W16506;
wire W16507;
wire W16508;
wire W16509;
wire W16510;
wire W16511;
wire W16512;
wire W16513;
wire W16514;
wire W16515;
wire W16516;
wire W16517;
wire W16518;
wire W16519;
wire W16520;
wire W16521;
wire W16522;
wire W16523;
wire W16524;
wire W16525;
wire W16526;
wire W16527;
wire W16528;
wire W16529;
wire W16530;
wire W16531;
wire W16532;
wire W16533;
wire W16534;
wire W16535;
wire W16536;
wire W16537;
wire W16538;
wire W16539;
wire W16540;
wire W16541;
wire W16542;
wire W16543;
wire W16544;
wire W16545;
wire W16546;
wire W16547;
wire W16548;
wire W16549;
wire W16550;
wire W16551;
wire W16552;
wire W16553;
wire W16554;
wire W16555;
wire W16556;
wire W16557;
wire W16558;
wire W16559;
wire W16560;
wire W16561;
wire W16562;
wire W16563;
wire W16564;
wire W16565;
wire W16566;
wire W16567;
wire W16568;
wire W16569;
wire W16570;
wire W16571;
wire W16572;
wire W16573;
wire W16574;
wire W16575;
wire W16576;
wire W16577;
wire W16578;
wire W16579;
wire W16580;
wire W16581;
wire W16582;
wire W16583;
wire W16584;
wire W16585;
wire W16586;
wire W16587;
wire W16588;
wire W16589;
wire W16590;
wire W16591;
wire W16592;
wire W16593;
wire W16594;
wire W16595;
wire W16596;
wire W16597;
wire W16598;
wire W16599;
wire W16600;
wire W16601;
wire W16602;
wire W16603;
wire W16604;
wire W16605;
wire W16606;
wire W16607;
wire W16608;
wire W16609;
wire W16610;
wire W16611;
wire W16612;
wire W16613;
wire W16614;
wire W16615;
wire W16616;
wire W16617;
wire W16618;
wire W16619;
wire W16620;
wire W16621;
wire W16622;
wire W16623;
wire W16624;
wire W16625;
wire W16626;
wire W16627;
wire W16628;
wire W16629;
wire W16630;
wire W16631;
wire W16632;
wire W16633;
wire W16634;
wire W16635;
wire W16636;
wire W16637;
wire W16638;
wire W16639;
wire W16640;
wire W16641;
wire W16642;
wire W16643;
wire W16644;
wire W16645;
wire W16646;
wire W16647;
wire W16648;
wire W16649;
wire W16650;
wire W16651;
wire W16652;
wire W16653;
wire W16654;
wire W16655;
wire W16656;
wire W16657;
wire W16658;
wire W16659;
wire W16660;
wire W16661;
wire W16662;
wire W16663;
wire W16664;
wire W16665;
wire W16666;
wire W16667;
wire W16668;
wire W16669;
wire W16670;
wire W16671;
wire W16672;
wire W16673;
wire W16674;
wire W16675;
wire W16676;
wire W16677;
wire W16678;
wire W16679;
wire W16680;
wire W16681;
wire W16682;
wire W16683;
wire W16684;
wire W16685;
wire W16686;
wire W16687;
wire W16688;
wire W16689;
wire W16690;
wire W16691;
wire W16692;
wire W16693;
wire W16694;
wire W16695;
wire W16696;
wire W16697;
wire W16698;
wire W16699;
wire W16700;
wire W16701;
wire W16702;
wire W16703;
wire W16704;
wire W16705;
wire W16706;
wire W16707;
wire W16708;
wire W16709;
wire W16710;
wire W16711;
wire W16712;
wire W16713;
wire W16714;
wire W16715;
wire W16716;
wire W16717;
wire W16718;
wire W16719;
wire W16720;
wire W16721;
wire W16722;
wire W16723;
wire W16724;
wire W16725;
wire W16726;
wire W16727;
wire W16728;
wire W16729;
wire W16730;
wire W16731;
wire W16732;
wire W16733;
wire W16734;
wire W16735;
wire W16736;
wire W16737;
wire W16738;
wire W16739;
wire W16740;
wire W16741;
wire W16742;
wire W16743;
wire W16744;
wire W16745;
wire W16746;
wire W16747;
wire W16748;
wire W16749;
wire W16750;
wire W16751;
wire W16752;
wire W16753;
wire W16754;
wire W16755;
wire W16756;
wire W16757;
wire W16758;
wire W16759;
wire W16760;
wire W16761;
wire W16762;
wire W16763;
wire W16764;
wire W16765;
wire W16766;
wire W16767;
wire W16768;
wire W16769;
wire W16770;
wire W16771;
wire W16772;
wire W16773;
wire W16774;
wire W16775;
wire W16776;
wire W16777;
wire W16778;
wire W16779;
wire W16780;
wire W16781;
wire W16782;
wire W16783;
wire W16784;
wire W16785;
wire W16786;
wire W16787;
wire W16788;
wire W16789;
wire W16790;
wire W16791;
wire W16792;
wire W16793;
wire W16794;
wire W16795;
wire W16796;
wire W16797;
wire W16798;
wire W16799;
wire W16800;
wire W16801;
wire W16802;
wire W16803;
wire W16804;
wire W16805;
wire W16806;
wire W16807;
wire W16808;
wire W16809;
wire W16810;
wire W16811;
wire W16812;
wire W16813;
wire W16814;
wire W16815;
wire W16816;
wire W16817;
wire W16818;
wire W16819;
wire W16820;
wire W16821;
wire W16822;
wire W16823;
wire W16824;
wire W16825;
wire W16826;
wire W16827;
wire W16828;
wire W16829;
wire W16830;
wire W16831;
wire W16832;
wire W16833;
wire W16834;
wire W16835;
wire W16836;
wire W16837;
wire W16838;
wire W16839;
wire W16840;
wire W16841;
wire W16842;
wire W16843;
wire W16844;
wire W16845;
wire W16846;
wire W16847;
wire W16848;
wire W16849;
wire W16850;
wire W16851;
wire W16852;
wire W16853;
wire W16854;
wire W16855;
wire W16856;
wire W16857;
wire W16858;
wire W16859;
wire W16860;
wire W16861;
wire W16862;
wire W16863;
wire W16864;
wire W16865;
wire W16866;
wire W16867;
wire W16868;
wire W16869;
wire W16870;
wire W16871;
wire W16872;
wire W16873;
wire W16874;
wire W16875;
wire W16876;
wire W16877;
wire W16878;
wire W16879;
wire W16880;
wire W16881;
wire W16882;
wire W16883;
wire W16884;
wire W16885;
wire W16886;
wire W16887;
wire W16888;
wire W16889;
wire W16890;
wire W16891;
wire W16892;
wire W16893;
wire W16894;
wire W16895;
wire W16896;
wire W16897;
wire W16898;
wire W16899;
wire W16900;
wire W16901;
wire W16902;
wire W16903;
wire W16904;
wire W16905;
wire W16906;
wire W16907;
wire W16908;
wire W16909;
wire W16910;
wire W16911;
wire W16912;
wire W16913;
wire W16914;
wire W16915;
wire W16916;
wire W16917;
wire W16918;
wire W16919;
wire W16920;
wire W16921;
wire W16922;
wire W16923;
wire W16924;
wire W16925;
wire W16926;
wire W16927;
wire W16928;
wire W16929;
wire W16930;
wire W16931;
wire W16932;
wire W16933;
wire W16934;
wire W16935;
wire W16936;
wire W16937;
wire W16938;
wire W16939;
wire W16940;
wire W16941;
wire W16942;
wire W16943;
wire W16944;
wire W16945;
wire W16946;
wire W16947;
wire W16948;
wire W16949;
wire W16950;
wire W16951;
wire W16952;
wire W16953;
wire W16954;
wire W16955;
wire W16956;
wire W16957;
wire W16958;
wire W16959;
wire W16960;
wire W16961;
wire W16962;
wire W16963;
wire W16964;
wire W16965;
wire W16966;
wire W16967;
wire W16968;
wire W16969;
wire W16970;
wire W16971;
wire W16972;
wire W16973;
wire W16974;
wire W16975;
wire W16976;
wire W16977;
wire W16978;
wire W16979;
wire W16980;
wire W16981;
wire W16982;
wire W16983;
wire W16984;
wire W16985;
wire W16986;
wire W16987;
wire W16988;
wire W16989;
wire W16990;
wire W16991;
wire W16992;
wire W16993;
wire W16994;
wire W16995;
wire W16996;
wire W16997;
wire W16998;
wire W16999;
wire W17000;
wire W17001;
wire W17002;
wire W17003;
wire W17004;
wire W17005;
wire W17006;
wire W17007;
wire W17008;
wire W17009;
wire W17010;
wire W17011;
wire W17012;
wire W17013;
wire W17014;
wire W17015;
wire W17016;
wire W17017;
wire W17018;
wire W17019;
wire W17020;
wire W17021;
wire W17022;
wire W17023;
wire W17024;
wire W17025;
wire W17026;
wire W17027;
wire W17028;
wire W17029;
wire W17030;
wire W17031;
wire W17032;
wire W17033;
wire W17034;
wire W17035;
wire W17036;
wire W17037;
wire W17038;
wire W17039;
wire W17040;
wire W17041;
wire W17042;
wire W17043;
wire W17044;
wire W17045;
wire W17046;
wire W17047;
wire W17048;
wire W17049;
wire W17050;
wire W17051;
wire W17052;
wire W17053;
wire W17054;
wire W17055;
wire W17056;
wire W17057;
wire W17058;
wire W17059;
wire W17060;
wire W17061;
wire W17062;
wire W17063;
wire W17064;
wire W17065;
wire W17066;
wire W17067;
wire W17068;
wire W17069;
wire W17070;
wire W17071;
wire W17072;
wire W17073;
wire W17074;
wire W17075;
wire W17076;
wire W17077;
wire W17078;
wire W17079;
wire W17080;
wire W17081;
wire W17082;
wire W17083;
wire W17084;
wire W17085;
wire W17086;
wire W17087;
wire W17088;
wire W17089;
wire W17090;
wire W17091;
wire W17092;
wire W17093;
wire W17094;
wire W17095;
wire W17096;
wire W17097;
wire W17098;
wire W17099;
wire W17100;
wire W17101;
wire W17102;
wire W17103;
wire W17104;
wire W17105;
wire W17106;
wire W17107;
wire W17108;
wire W17109;
wire W17110;
wire W17111;
wire W17112;
wire W17113;
wire W17114;
wire W17115;
wire W17116;
wire W17117;
wire W17118;
wire W17119;
wire W17120;
wire W17121;
wire W17122;
wire W17123;
wire W17124;
wire W17125;
wire W17126;
wire W17127;
wire W17128;
wire W17129;
wire W17130;
wire W17131;
wire W17132;
wire W17133;
wire W17134;
wire W17135;
wire W17136;
wire W17137;
wire W17138;
wire W17139;
wire W17140;
wire W17141;
wire W17142;
wire W17143;
wire W17144;
wire W17145;
wire W17146;
wire W17147;
wire W17148;
wire W17149;
wire W17150;
wire W17151;
wire W17152;
wire W17153;
wire W17154;
wire W17155;
wire W17156;
wire W17157;
wire W17158;
wire W17159;
wire W17160;
wire W17161;
wire W17162;
wire W17163;
wire W17164;
wire W17165;
wire W17166;
wire W17167;
wire W17168;
wire W17169;
wire W17170;
wire W17171;
wire W17172;
wire W17173;
wire W17174;
wire W17175;
wire W17176;
wire W17177;
wire W17178;
wire W17179;
wire W17180;
wire W17181;
wire W17182;
wire W17183;
wire W17184;
wire W17185;
wire W17186;
wire W17187;
wire W17188;
wire W17189;
wire W17190;
wire W17191;
wire W17192;
wire W17193;
wire W17194;
wire W17195;
wire W17196;
wire W17197;
wire W17198;
wire W17199;
wire W17200;
wire W17201;
wire W17202;
wire W17203;
wire W17204;
wire W17205;
wire W17206;
wire W17207;
wire W17208;
wire W17209;
wire W17210;
wire W17211;
wire W17212;
wire W17213;
wire W17214;
wire W17215;
wire W17216;
wire W17217;
wire W17218;
wire W17219;
wire W17220;
wire W17221;
wire W17222;
wire W17223;
wire W17224;
wire W17225;
wire W17226;
wire W17227;
wire W17228;
wire W17229;
wire W17230;
wire W17231;
wire W17232;
wire W17233;
wire W17234;
wire W17235;
wire W17236;
wire W17237;
wire W17238;
wire W17239;
wire W17240;
wire W17241;
wire W17242;
wire W17243;
wire W17244;
wire W17245;
wire W17246;
wire W17247;
wire W17248;
wire W17249;
wire W17250;
wire W17251;
wire W17252;
wire W17253;
wire W17254;
wire W17255;
wire W17256;
wire W17257;
wire W17258;
wire W17259;
wire W17260;
wire W17261;
wire W17262;
wire W17263;
wire W17264;
wire W17265;
wire W17266;
wire W17267;
wire W17268;
wire W17269;
wire W17270;
wire W17271;
wire W17272;
wire W17273;
wire W17274;
wire W17275;
wire W17276;
wire W17277;
wire W17278;
wire W17279;
wire W17280;
wire W17281;
wire W17282;
wire W17283;
wire W17284;
wire W17285;
wire W17286;
wire W17287;
wire W17288;
wire W17289;
wire W17290;
wire W17291;
wire W17292;
wire W17293;
wire W17294;
wire W17295;
wire W17296;
wire W17297;
wire W17298;
wire W17299;
wire W17300;
wire W17301;
wire W17302;
wire W17303;
wire W17304;
wire W17305;
wire W17306;
wire W17307;
wire W17308;
wire W17309;
wire W17310;
wire W17311;
wire W17312;
wire W17313;
wire W17314;
wire W17315;
wire W17316;
wire W17317;
wire W17318;
wire W17319;
wire W17320;
wire W17321;
wire W17322;
wire W17323;
wire W17324;
wire W17325;
wire W17326;
wire W17327;
wire W17328;
wire W17329;
wire W17330;
wire W17331;
wire W17332;
wire W17333;
wire W17334;
wire W17335;
wire W17336;
wire W17337;
wire W17338;
wire W17339;
wire W17340;
wire W17341;
wire W17342;
wire W17343;
wire W17344;
wire W17345;
wire W17346;
wire W17347;
wire W17348;
wire W17349;
wire W17350;
wire W17351;
wire W17352;
wire W17353;
wire W17354;
wire W17355;
wire W17356;
wire W17357;
wire W17358;
wire W17359;
wire W17360;
wire W17361;
wire W17362;
wire W17363;
wire W17364;
wire W17365;
wire W17366;
wire W17367;
wire W17368;
wire W17369;
wire W17370;
wire W17371;
wire W17372;
wire W17373;
wire W17374;
wire W17375;
wire W17376;
wire W17377;
wire W17378;
wire W17379;
wire W17380;
wire W17381;
wire W17382;
wire W17383;
wire W17384;
wire W17385;
wire W17386;
wire W17387;
wire W17388;
wire W17389;
wire W17390;
wire W17391;
wire W17392;
wire W17393;
wire W17394;
wire W17395;
wire W17396;
wire W17397;
wire W17398;
wire W17399;
wire W17400;
wire W17401;
wire W17402;
wire W17403;
wire W17404;
wire W17405;
wire W17406;
wire W17407;
wire W17408;
wire W17409;
wire W17410;
wire W17411;
wire W17412;
wire W17413;
wire W17414;
wire W17415;
wire W17416;
wire W17417;
wire W17418;
wire W17419;
wire W17420;
wire W17421;
wire W17422;
wire W17423;
wire W17424;
wire W17425;
wire W17426;
wire W17427;
wire W17428;
wire W17429;
wire W17430;
wire W17431;
wire W17432;
wire W17433;
wire W17434;
wire W17435;
wire W17436;
wire W17437;
wire W17438;
wire W17439;
wire W17440;
wire W17441;
wire W17442;
wire W17443;
wire W17444;
wire W17445;
wire W17446;
wire W17447;
wire W17448;
wire W17449;
wire W17450;
wire W17451;
wire W17452;
wire W17453;
wire W17454;
wire W17455;
wire W17456;
wire W17457;
wire W17458;
wire W17459;
wire W17460;
wire W17461;
wire W17462;
wire W17463;
wire W17464;
wire W17465;
wire W17466;
wire W17467;
wire W17468;
wire W17469;
wire W17470;
wire W17471;
wire W17472;
wire W17473;
wire W17474;
wire W17475;
wire W17476;
wire W17477;
wire W17478;
wire W17479;
wire W17480;
wire W17481;
wire W17482;
wire W17483;
wire W17484;
wire W17485;
wire W17486;
wire W17487;
wire W17488;
wire W17489;
wire W17490;
wire W17491;
wire W17492;
wire W17493;
wire W17494;
wire W17495;
wire W17496;
wire W17497;
wire W17498;
wire W17499;
wire W17500;
wire W17501;
wire W17502;
wire W17503;
wire W17504;
wire W17505;
wire W17506;
wire W17507;
wire W17508;
wire W17509;
wire W17510;
wire W17511;
wire W17512;
wire W17513;
wire W17514;
wire W17515;
wire W17516;
wire W17517;
wire W17518;
wire W17519;
wire W17520;
wire W17521;
wire W17522;
wire W17523;
wire W17524;
wire W17525;
wire W17526;
wire W17527;
wire W17528;
wire W17529;
wire W17530;
wire W17531;
wire W17532;
wire W17533;
wire W17534;
wire W17535;
wire W17536;
wire W17537;
wire W17538;
wire W17539;
wire W17540;
wire W17541;
wire W17542;
wire W17543;
wire W17544;
wire W17545;
wire W17546;
wire W17547;
wire W17548;
wire W17549;
wire W17550;
wire W17551;
wire W17552;
wire W17553;
wire W17554;
wire W17555;
wire W17556;
wire W17557;
wire W17558;
wire W17559;
wire W17560;
wire W17561;
wire W17562;
wire W17563;
wire W17564;
wire W17565;
wire W17566;
wire W17567;
wire W17568;
wire W17569;
wire W17570;
wire W17571;
wire W17572;
wire W17573;
wire W17574;
wire W17575;
wire W17576;
wire W17577;
wire W17578;
wire W17579;
wire W17580;
wire W17581;
wire W17582;
wire W17583;
wire W17584;
wire W17585;
wire W17586;
wire W17587;
wire W17588;
wire W17589;
wire W17590;
wire W17591;
wire W17592;
wire W17593;
wire W17594;
wire W17595;
wire W17596;
wire W17597;
wire W17598;
wire W17599;
wire W17600;
wire W17601;
wire W17602;
wire W17603;
wire W17604;
wire W17605;
wire W17606;
wire W17607;
wire W17608;
wire W17609;
wire W17610;
wire W17611;
wire W17612;
wire W17613;
wire W17614;
wire W17615;
wire W17616;
wire W17617;
wire W17618;
wire W17619;
wire W17620;
wire W17621;
wire W17622;
wire W17623;
wire W17624;
wire W17625;
wire W17626;
wire W17627;
wire W17628;
wire W17629;
wire W17630;
wire W17631;
wire W17632;
wire W17633;
wire W17634;
wire W17635;
wire W17636;
wire W17637;
wire W17638;
wire W17639;
wire W17640;
wire W17641;
wire W17642;
wire W17643;
wire W17644;
wire W17645;
wire W17646;
wire W17647;
wire W17648;
wire W17649;
wire W17650;
wire W17651;
wire W17652;
wire W17653;
wire W17654;
wire W17655;
wire W17656;
wire W17657;
wire W17658;
wire W17659;
wire W17660;
wire W17661;
wire W17662;
wire W17663;
wire W17664;
wire W17665;
wire W17666;
wire W17667;
wire W17668;
wire W17669;
wire W17670;
wire W17671;
wire W17672;
wire W17673;
wire W17674;
wire W17675;
wire W17676;
wire W17677;
wire W17678;
wire W17679;
wire W17680;
wire W17681;
wire W17682;
wire W17683;
wire W17684;
wire W17685;
wire W17686;
wire W17687;
wire W17688;
wire W17689;
wire W17690;
wire W17691;
wire W17692;
wire W17693;
wire W17694;
wire W17695;
wire W17696;
wire W17697;
wire W17698;
wire W17699;
wire W17700;
wire W17701;
wire W17702;
wire W17703;
wire W17704;
wire W17705;
wire W17706;
wire W17707;
wire W17708;
wire W17709;
wire W17710;
wire W17711;
wire W17712;
wire W17713;
wire W17714;
wire W17715;
wire W17716;
wire W17717;
wire W17718;
wire W17719;
wire W17720;
wire W17721;
wire W17722;
wire W17723;
wire W17724;
wire W17725;
wire W17726;
wire W17727;
wire W17728;
wire W17729;
wire W17730;
wire W17731;
wire W17732;
wire W17733;
wire W17734;
wire W17735;
wire W17736;
wire W17737;
wire W17738;
wire W17739;
wire W17740;
wire W17741;
wire W17742;
wire W17743;
wire W17744;
wire W17745;
wire W17746;
wire W17747;
wire W17748;
wire W17749;
wire W17750;
wire W17751;
wire W17752;
wire W17753;
wire W17754;
wire W17755;
wire W17756;
wire W17757;
wire W17758;
wire W17759;
wire W17760;
wire W17761;
wire W17762;
wire W17763;
wire W17764;
wire W17765;
wire W17766;
wire W17767;
wire W17768;
wire W17769;
wire W17770;
wire W17771;
wire W17772;
wire W17773;
wire W17774;
wire W17775;
wire W17776;
wire W17777;
wire W17778;
wire W17779;
wire W17780;
wire W17781;
wire W17782;
wire W17783;
wire W17784;
wire W17785;
wire W17786;
wire W17787;
wire W17788;
wire W17789;
wire W17790;
wire W17791;
wire W17792;
wire W17793;
wire W17794;
wire W17795;
wire W17796;
wire W17797;
wire W17798;
wire W17799;
wire W17800;
wire W17801;
wire W17802;
wire W17803;
wire W17804;
wire W17805;
wire W17806;
wire W17807;
wire W17808;
wire W17809;
wire W17810;
wire W17811;
wire W17812;
wire W17813;
wire W17814;
wire W17815;
wire W17816;
wire W17817;
wire W17818;
wire W17819;
wire W17820;
wire W17821;
wire W17822;
wire W17823;
wire W17824;
wire W17825;
wire W17826;
wire W17827;
wire W17828;
wire W17829;
wire W17830;
wire W17831;
wire W17832;
wire W17833;
wire W17834;
wire W17835;
wire W17836;
wire W17837;
wire W17838;
wire W17839;
wire W17840;
wire W17841;
wire W17842;
wire W17843;
wire W17844;
wire W17845;
wire W17846;
wire W17847;
wire W17848;
wire W17849;
wire W17850;
wire W17851;
wire W17852;
wire W17853;
wire W17854;
wire W17855;
wire W17856;
wire W17857;
wire W17858;
wire W17859;
wire W17860;
wire W17861;
wire W17862;
wire W17863;
wire W17864;
wire W17865;
wire W17866;
wire W17867;
wire W17868;
wire W17869;
wire W17870;
wire W17871;
wire W17872;
wire W17873;
wire W17874;
wire W17875;
wire W17876;
wire W17877;
wire W17878;
wire W17879;
wire W17880;
wire W17881;
wire W17882;
wire W17883;
wire W17884;
wire W17885;
wire W17886;
wire W17887;
wire W17888;
wire W17889;
wire W17890;
wire W17891;
wire W17892;
wire W17893;
wire W17894;
wire W17895;
wire W17896;
wire W17897;
wire W17898;
wire W17899;
wire W17900;
wire W17901;
wire W17902;
wire W17903;
wire W17904;
wire W17905;
wire W17906;
wire W17907;
wire W17908;
wire W17909;
wire W17910;
wire W17911;
wire W17912;
wire W17913;
wire W17914;
wire W17915;
wire W17916;
wire W17917;
wire W17918;
wire W17919;
wire W17920;
wire W17921;
wire W17922;
wire W17923;
wire W17924;
wire W17925;
wire W17926;
wire W17927;
wire W17928;
wire W17929;
wire W17930;
wire W17931;
wire W17932;
wire W17933;
wire W17934;
wire W17935;
wire W17936;
wire W17937;
wire W17938;
wire W17939;
wire W17940;
wire W17941;
wire W17942;
wire W17943;
wire W17944;
wire W17945;
wire W17946;
wire W17947;
wire W17948;
wire W17949;
wire W17950;
wire W17951;
wire W17952;
wire W17953;
wire W17954;
wire W17955;
wire W17956;
wire W17957;
wire W17958;
wire W17959;
wire W17960;
wire W17961;
wire W17962;
wire W17963;
wire W17964;
wire W17965;
wire W17966;
wire W17967;
wire W17968;
wire W17969;
wire W17970;
wire W17971;
wire W17972;
wire W17973;
wire W17974;
wire W17975;
wire W17976;
wire W17977;
wire W17978;
wire W17979;
wire W17980;
wire W17981;
wire W17982;
wire W17983;
wire W17984;
wire W17985;
wire W17986;
wire W17987;
wire W17988;
wire W17989;
wire W17990;
wire W17991;
wire W17992;
wire W17993;
wire W17994;
wire W17995;
wire W17996;
wire W17997;
wire W17998;
wire W17999;
wire W18000;
wire W18001;
wire W18002;
wire W18003;
wire W18004;
wire W18005;
wire W18006;
wire W18007;
wire W18008;
wire W18009;
wire W18010;
wire W18011;
wire W18012;
wire W18013;
wire W18014;
wire W18015;
wire W18016;
wire W18017;
wire W18018;
wire W18019;
wire W18020;
wire W18021;
wire W18022;
wire W18023;
wire W18024;
wire W18025;
wire W18026;
wire W18027;
wire W18028;
wire W18029;
wire W18030;
wire W18031;
wire W18032;
wire W18033;
wire W18034;
wire W18035;
wire W18036;
wire W18037;
wire W18038;
wire W18039;
wire W18040;
wire W18041;
wire W18042;
wire W18043;
wire W18044;
wire W18045;
wire W18046;
wire W18047;
wire W18048;
wire W18049;
wire W18050;
wire W18051;
wire W18052;
wire W18053;
wire W18054;
wire W18055;
wire W18056;
wire W18057;
wire W18058;
wire W18059;
wire W18060;
wire W18061;
wire W18062;
wire W18063;
wire W18064;
wire W18065;
wire W18066;
wire W18067;
wire W18068;
wire W18069;
wire W18070;
wire W18071;
wire W18072;
wire W18073;
wire W18074;
wire W18075;
wire W18076;
wire W18077;
wire W18078;
wire W18079;
wire W18080;
wire W18081;
wire W18082;
wire W18083;
wire W18084;
wire W18085;
wire W18086;
wire W18087;
wire W18088;
wire W18089;
wire W18090;
wire W18091;
wire W18092;
wire W18093;
wire W18094;
wire W18095;
wire W18096;
wire W18097;
wire W18098;
wire W18099;
wire W18100;
wire W18101;
wire W18102;
wire W18103;
wire W18104;
wire W18105;
wire W18106;
wire W18107;
wire W18108;
wire W18109;
wire W18110;
wire W18111;
wire W18112;
wire W18113;
wire W18114;
wire W18115;
wire W18116;
wire W18117;
wire W18118;
wire W18119;
wire W18120;
wire W18121;
wire W18122;
wire W18123;
wire W18124;
wire W18125;
wire W18126;
wire W18127;
wire W18128;
wire W18129;
wire W18130;
wire W18131;
wire W18132;
wire W18133;
wire W18134;
wire W18135;
wire W18136;
wire W18137;
wire W18138;
wire W18139;
wire W18140;
wire W18141;
wire W18142;
wire W18143;
wire W18144;
wire W18145;
wire W18146;
wire W18147;
wire W18148;
wire W18149;
wire W18150;
wire W18151;
wire W18152;
wire W18153;
wire W18154;
wire W18155;
wire W18156;
wire W18157;
wire W18158;
wire W18159;
wire W18160;
wire W18161;
wire W18162;
wire W18163;
wire W18164;
wire W18165;
wire W18166;
wire W18167;
wire W18168;
wire W18169;
wire W18170;
wire W18171;
wire W18172;
wire W18173;
wire W18174;
wire W18175;
wire W18176;
wire W18177;
wire W18178;
wire W18179;
wire W18180;
wire W18181;
wire W18182;
wire W18183;
wire W18184;
wire W18185;
wire W18186;
wire W18187;
wire W18188;
wire W18189;
wire W18190;
wire W18191;
wire W18192;
wire W18193;
wire W18194;
wire W18195;
wire W18196;
wire W18197;
wire W18198;
wire W18199;
wire W18200;
wire W18201;
wire W18202;
wire W18203;
wire W18204;
wire W18205;
wire W18206;
wire W18207;
wire W18208;
wire W18209;
wire W18210;
wire W18211;
wire W18212;
wire W18213;
wire W18214;
wire W18215;
wire W18216;
wire W18217;
wire W18218;
wire W18219;
wire W18220;
wire W18221;
wire W18222;
wire W18223;
wire W18224;
wire W18225;
wire W18226;
wire W18227;
wire W18228;
wire W18229;
wire W18230;
wire W18231;
wire W18232;
wire W18233;
wire W18234;
wire W18235;
wire W18236;
wire W18237;
wire W18238;
wire W18239;
wire W18240;
wire W18241;
wire W18242;
wire W18243;
wire W18244;
wire W18245;
wire W18246;
wire W18247;
wire W18248;
wire W18249;
wire W18250;
wire W18251;
wire W18252;
wire W18253;
wire W18254;
wire W18255;
wire W18256;
wire W18257;
wire W18258;
wire W18259;
wire W18260;
wire W18261;
wire W18262;
wire W18263;
wire W18264;
wire W18265;
wire W18266;
wire W18267;
wire W18268;
wire W18269;
wire W18270;
wire W18271;
wire W18272;
wire W18273;
wire W18274;
wire W18275;
wire W18276;
wire W18277;
wire W18278;
wire W18279;
wire W18280;
wire W18281;
wire W18282;
wire W18283;
wire W18284;
wire W18285;
wire W18286;
wire W18287;
wire W18288;
wire W18289;
wire W18290;
wire W18291;
wire W18292;
wire W18293;
wire W18294;
wire W18295;
wire W18296;
wire W18297;
wire W18298;
wire W18299;
wire W18300;
wire W18301;
wire W18302;
wire W18303;
wire W18304;
wire W18305;
wire W18306;
wire W18307;
wire W18308;
wire W18309;
wire W18310;
wire W18311;
wire W18312;
wire W18313;
wire W18314;
wire W18315;
wire W18316;
wire W18317;
wire W18318;
wire W18319;
wire W18320;
wire W18321;
wire W18322;
wire W18323;
wire W18324;
wire W18325;
wire W18326;
wire W18327;
wire W18328;
wire W18329;
wire W18330;
wire W18331;
wire W18332;
wire W18333;
wire W18334;
wire W18335;
wire W18336;
wire W18337;
wire W18338;
wire W18339;
wire W18340;
wire W18341;
wire W18342;
wire W18343;
wire W18344;
wire W18345;
wire W18346;
wire W18347;
wire W18348;
wire W18349;
wire W18350;
wire W18351;
wire W18352;
wire W18353;
wire W18354;
wire W18355;
wire W18356;
wire W18357;
wire W18358;
wire W18359;
wire W18360;
wire W18361;
wire W18362;
wire W18363;
wire W18364;
wire W18365;
wire W18366;
wire W18367;
wire W18368;
wire W18369;
wire W18370;
wire W18371;
wire W18372;
wire W18373;
wire W18374;
wire W18375;
wire W18376;
wire W18377;
wire W18378;
wire W18379;
wire W18380;
wire W18381;
wire W18382;
wire W18383;
wire W18384;
wire W18385;
wire W18386;
wire W18387;
wire W18388;
wire W18389;
wire W18390;
wire W18391;
wire W18392;
wire W18393;
wire W18394;
wire W18395;
wire W18396;
wire W18397;
wire W18398;
wire W18399;
wire W18400;
wire W18401;
wire W18402;
wire W18403;
wire W18404;
wire W18405;
wire W18406;
wire W18407;
wire W18408;
wire W18409;
wire W18410;
wire W18411;
wire W18412;
wire W18413;
wire W18414;
wire W18415;
wire W18416;
wire W18417;
wire W18418;
wire W18419;
wire W18420;
wire W18421;
wire W18422;
wire W18423;
wire W18424;
wire W18425;
wire W18426;
wire W18427;
wire W18428;
wire W18429;
wire W18430;
wire W18431;
wire W18432;
wire W18433;
wire W18434;
wire W18435;
wire W18436;
wire W18437;
wire W18438;
wire W18439;
wire W18440;
wire W18441;
wire W18442;
wire W18443;
wire W18444;
wire W18445;
wire W18446;
wire W18447;
wire W18448;
wire W18449;
wire W18450;
wire W18451;
wire W18452;
wire W18453;
wire W18454;
wire W18455;
wire W18456;
wire W18457;
wire W18458;
wire W18459;
wire W18460;
wire W18461;
wire W18462;
wire W18463;
wire W18464;
wire W18465;
wire W18466;
wire W18467;
wire W18468;
wire W18469;
wire W18470;
wire W18471;
wire W18472;
wire W18473;
wire W18474;
wire W18475;
wire W18476;
wire W18477;
wire W18478;
wire W18479;
wire W18480;
wire W18481;
wire W18482;
wire W18483;
wire W18484;
wire W18485;
wire W18486;
wire W18487;
wire W18488;
wire W18489;
wire W18490;
wire W18491;
wire W18492;
wire W18493;
wire W18494;
wire W18495;
wire W18496;
wire W18497;
wire W18498;
wire W18499;
wire W18500;
wire W18501;
wire W18502;
wire W18503;
wire W18504;
wire W18505;
wire W18506;
wire W18507;
wire W18508;
wire W18509;
wire W18510;
wire W18511;
wire W18512;
wire W18513;
wire W18514;
wire W18515;
wire W18516;
wire W18517;
wire W18518;
wire W18519;
wire W18520;
wire W18521;
wire W18522;
wire W18523;
wire W18524;
wire W18525;
wire W18526;
wire W18527;
wire W18528;
wire W18529;
wire W18530;
wire W18531;
wire W18532;
wire W18533;
wire W18534;
wire W18535;
wire W18536;
wire W18537;
wire W18538;
wire W18539;
wire W18540;
wire W18541;
wire W18542;
wire W18543;
wire W18544;
wire W18545;
wire W18546;
wire W18547;
wire W18548;
wire W18549;
wire W18550;
wire W18551;
wire W18552;
wire W18553;
wire W18554;
wire W18555;
wire W18556;
wire W18557;
wire W18558;
wire W18559;
wire W18560;
wire W18561;
wire W18562;
wire W18563;
wire W18564;
wire W18565;
wire W18566;
wire W18567;
wire W18568;
wire W18569;
wire W18570;
wire W18571;
wire W18572;
wire W18573;
wire W18574;
wire W18575;
wire W18576;
wire W18577;
wire W18578;
wire W18579;
wire W18580;
wire W18581;
wire W18582;
wire W18583;
wire W18584;
wire W18585;
wire W18586;
wire W18587;
wire W18588;
wire W18589;
wire W18590;
wire W18591;
wire W18592;
wire W18593;
wire W18594;
wire W18595;
wire W18596;
wire W18597;
wire W18598;
wire W18599;
wire W18600;
wire W18601;
wire W18602;
wire W18603;
wire W18604;
wire W18605;
wire W18606;
wire W18607;
wire W18608;
wire W18609;
wire W18610;
wire W18611;
wire W18612;
wire W18613;
wire W18614;
wire W18615;
wire W18616;
wire W18617;
wire W18618;
wire W18619;
wire W18620;
wire W18621;
wire W18622;
wire W18623;
wire W18624;
wire W18625;
wire W18626;
wire W18627;
wire W18628;
wire W18629;
wire W18630;
wire W18631;
wire W18632;
wire W18633;
wire W18634;
wire W18635;
wire W18636;
wire W18637;
wire W18638;
wire W18639;
wire W18640;
wire W18641;
wire W18642;
wire W18643;
wire W18644;
wire W18645;
wire W18646;
wire W18647;
wire W18648;
wire W18649;
wire W18650;
wire W18651;
wire W18652;
wire W18653;
wire W18654;
wire W18655;
wire W18656;
wire W18657;
wire W18658;
wire W18659;
wire W18660;
wire W18661;
wire W18662;
wire W18663;
wire W18664;
wire W18665;
wire W18666;
wire W18667;
wire W18668;
wire W18669;
wire W18670;
wire W18671;
wire W18672;
wire W18673;
wire W18674;
wire W18675;
wire W18676;
wire W18677;
wire W18678;
wire W18679;
wire W18680;
wire W18681;
wire W18682;
wire W18683;
wire W18684;
wire W18685;
wire W18686;
wire W18687;
wire W18688;
wire W18689;
wire W18690;
wire W18691;
wire W18692;
wire W18693;
wire W18694;
wire W18695;
wire W18696;
wire W18697;
wire W18698;
wire W18699;
wire W18700;
wire W18701;
wire W18702;
wire W18703;
wire W18704;
wire W18705;
wire W18706;
wire W18707;
wire W18708;
wire W18709;
wire W18710;
wire W18711;
wire W18712;
wire W18713;
wire W18714;
wire W18715;
wire W18716;
wire W18717;
wire W18718;
wire W18719;
wire W18720;
wire W18721;
wire W18722;
wire W18723;
wire W18724;
wire W18725;
wire W18726;
wire W18727;
wire W18728;
wire W18729;
wire W18730;
wire W18731;
wire W18732;
wire W18733;
wire W18734;
wire W18735;
wire W18736;
wire W18737;
wire W18738;
wire W18739;
wire W18740;
wire W18741;
wire W18742;
wire W18743;
wire W18744;
wire W18745;
wire W18746;
wire W18747;
wire W18748;
wire W18749;
wire W18750;
wire W18751;
wire W18752;
wire W18753;
wire W18754;
wire W18755;
wire W18756;
wire W18757;
wire W18758;
wire W18759;
wire W18760;
wire W18761;
wire W18762;
wire W18763;
wire W18764;
wire W18765;
wire W18766;
wire W18767;
wire W18768;
wire W18769;
wire W18770;
wire W18771;
wire W18772;
wire W18773;
wire W18774;
wire W18775;
wire W18776;
wire W18777;
wire W18778;
wire W18779;
wire W18780;
wire W18781;
wire W18782;
wire W18783;
wire W18784;
wire W18785;
wire W18786;
wire W18787;
wire W18788;
wire W18789;
wire W18790;
wire W18791;
wire W18792;
wire W18793;
wire W18794;
wire W18795;
wire W18796;
wire W18797;
wire W18798;
wire W18799;
wire W18800;
wire W18801;
wire W18802;
wire W18803;
wire W18804;
wire W18805;
wire W18806;
wire W18807;
wire W18808;
wire W18809;
wire W18810;
wire W18811;
wire W18812;
wire W18813;
wire W18814;
wire W18815;
wire W18816;
wire W18817;
wire W18818;
wire W18819;
wire W18820;
wire W18821;
wire W18822;
wire W18823;
wire W18824;
wire W18825;
wire W18826;
wire W18827;
wire W18828;
wire W18829;
wire W18830;
wire W18831;
wire W18832;
wire W18833;
wire W18834;
wire W18835;
wire W18836;
wire W18837;
wire W18838;
wire W18839;
wire W18840;
wire W18841;
wire W18842;
wire W18843;
wire W18844;
wire W18845;
wire W18846;
wire W18847;
wire W18848;
wire W18849;
wire W18850;
wire W18851;
wire W18852;
wire W18853;
wire W18854;
wire W18855;
wire W18856;
wire W18857;
wire W18858;
wire W18859;
wire W18860;
wire W18861;
wire W18862;
wire W18863;
wire W18864;
wire W18865;
wire W18866;
wire W18867;
wire W18868;
wire W18869;
wire W18870;
wire W18871;
wire W18872;
wire W18873;
wire W18874;
wire W18875;
wire W18876;
wire W18877;
wire W18878;
wire W18879;
wire W18880;
wire W18881;
wire W18882;
wire W18883;
wire W18884;
wire W18885;
wire W18886;
wire W18887;
wire W18888;
wire W18889;
wire W18890;
wire W18891;
wire W18892;
wire W18893;
wire W18894;
wire W18895;
wire W18896;
wire W18897;
wire W18898;
wire W18899;
wire W18900;
wire W18901;
wire W18902;
wire W18903;
wire W18904;
wire W18905;
wire W18906;
wire W18907;
wire W18908;
wire W18909;
wire W18910;
wire W18911;
wire W18912;
wire W18913;
wire W18914;
wire W18915;
wire W18916;
wire W18917;
wire W18918;
wire W18919;
wire W18920;
wire W18921;
wire W18922;
wire W18923;
wire W18924;
wire W18925;
wire W18926;
wire W18927;
wire W18928;
wire W18929;
wire W18930;
wire W18931;
wire W18932;
wire W18933;
wire W18934;
wire W18935;
wire W18936;
wire W18937;
wire W18938;
wire W18939;
wire W18940;
wire W18941;
wire W18942;
wire W18943;
wire W18944;
wire W18945;
wire W18946;
wire W18947;
wire W18948;
wire W18949;
wire W18950;
wire W18951;
wire W18952;
wire W18953;
wire W18954;
wire W18955;
wire W18956;
wire W18957;
wire W18958;
wire W18959;
wire W18960;
wire W18961;
wire W18962;
wire W18963;
wire W18964;
wire W18965;
wire W18966;
wire W18967;
wire W18968;
wire W18969;
wire W18970;
wire W18971;
wire W18972;
wire W18973;
wire W18974;
wire W18975;
wire W18976;
wire W18977;
wire W18978;
wire W18979;
wire W18980;
wire W18981;
wire W18982;
wire W18983;
wire W18984;
wire W18985;
wire W18986;
wire W18987;
wire W18988;
wire W18989;
wire W18990;
wire W18991;
wire W18992;
wire W18993;
wire W18994;
wire W18995;
wire W18996;
wire W18997;
wire W18998;
wire W18999;
wire W19000;
wire W19001;
wire W19002;
wire W19003;
wire W19004;
wire W19005;
wire W19006;
wire W19007;
wire W19008;
wire W19009;
wire W19010;
wire W19011;
wire W19012;
wire W19013;
wire W19014;
wire W19015;
wire W19016;
wire W19017;
wire W19018;
wire W19019;
wire W19020;
wire W19021;
wire W19022;
wire W19023;
wire W19024;
wire W19025;
wire W19026;
wire W19027;
wire W19028;
wire W19029;
wire W19030;
wire W19031;
wire W19032;
wire W19033;
wire W19034;
wire W19035;
wire W19036;
wire W19037;
wire W19038;
wire W19039;
wire W19040;
wire W19041;
wire W19042;
wire W19043;
wire W19044;
wire W19045;
wire W19046;
wire W19047;
wire W19048;
wire W19049;
wire W19050;
wire W19051;
wire W19052;
wire W19053;
wire W19054;
wire W19055;
wire W19056;
wire W19057;
wire W19058;
wire W19059;
wire W19060;
wire W19061;
wire W19062;
wire W19063;
wire W19064;
wire W19065;
wire W19066;
wire W19067;
wire W19068;
wire W19069;
wire W19070;
wire W19071;
wire W19072;
wire W19073;
wire W19074;
wire W19075;
wire W19076;
wire W19077;
wire W19078;
wire W19079;
wire W19080;
wire W19081;
wire W19082;
wire W19083;
wire W19084;
wire W19085;
wire W19086;
wire W19087;
wire W19088;
wire W19089;
wire W19090;
wire W19091;
wire W19092;
wire W19093;
wire W19094;
wire W19095;
wire W19096;
wire W19097;
wire W19098;
wire W19099;
wire W19100;
wire W19101;
wire W19102;
wire W19103;
wire W19104;
wire W19105;
wire W19106;
wire W19107;
wire W19108;
wire W19109;
wire W19110;
wire W19111;
wire W19112;
wire W19113;
wire W19114;
wire W19115;
wire W19116;
wire W19117;
wire W19118;
wire W19119;
wire W19120;
wire W19121;
wire W19122;
wire W19123;
wire W19124;
wire W19125;
wire W19126;
wire W19127;
wire W19128;
wire W19129;
wire W19130;
wire W19131;
wire W19132;
wire W19133;
wire W19134;
wire W19135;
wire W19136;
wire W19137;
wire W19138;
wire W19139;
wire W19140;
wire W19141;
wire W19142;
wire W19143;
wire W19144;
wire W19145;
wire W19146;
wire W19147;
wire W19148;
wire W19149;
wire W19150;
wire W19151;
wire W19152;
wire W19153;
wire W19154;
wire W19155;
wire W19156;
wire W19157;
wire W19158;
wire W19159;
wire W19160;
wire W19161;
wire W19162;
wire W19163;
wire W19164;
wire W19165;
wire W19166;
wire W19167;
wire W19168;
wire W19169;
wire W19170;
wire W19171;
wire W19172;
wire W19173;
wire W19174;
wire W19175;
wire W19176;
wire W19177;
wire W19178;
wire W19179;
wire W19180;
wire W19181;
wire W19182;
wire W19183;
wire W19184;
wire W19185;
wire W19186;
wire W19187;
wire W19188;
wire W19189;
wire W19190;
wire W19191;
wire W19192;
wire W19193;
wire W19194;
wire W19195;
wire W19196;
wire W19197;
wire W19198;
wire W19199;
wire W19200;
wire W19201;
wire W19202;
wire W19203;
wire W19204;
wire W19205;
wire W19206;
wire W19207;
wire W19208;
wire W19209;
wire W19210;
wire W19211;
wire W19212;
wire W19213;
wire W19214;
wire W19215;
wire W19216;
wire W19217;
wire W19218;
wire W19219;
wire W19220;
wire W19221;
wire W19222;
wire W19223;
wire W19224;
wire W19225;
wire W19226;
wire W19227;
wire W19228;
wire W19229;
wire W19230;
wire W19231;
wire W19232;
wire W19233;
wire W19234;
wire W19235;
wire W19236;
wire W19237;
wire W19238;
wire W19239;
wire W19240;
wire W19241;
wire W19242;
wire W19243;
wire W19244;
wire W19245;
wire W19246;
wire W19247;
wire W19248;
wire W19249;
wire W19250;
wire W19251;
wire W19252;
wire W19253;
wire W19254;
wire W19255;
wire W19256;
wire W19257;
wire W19258;
wire W19259;
wire W19260;
wire W19261;
wire W19262;
wire W19263;
wire W19264;
wire W19265;
wire W19266;
wire W19267;
wire W19268;
wire W19269;
wire W19270;
wire W19271;
wire W19272;
wire W19273;
wire W19274;
wire W19275;
wire W19276;
wire W19277;
wire W19278;
wire W19279;
wire W19280;
wire W19281;
wire W19282;
wire W19283;
wire W19284;
wire W19285;
wire W19286;
wire W19287;
wire W19288;
wire W19289;
wire W19290;
wire W19291;
wire W19292;
wire W19293;
wire W19294;
wire W19295;
wire W19296;
wire W19297;
wire W19298;
wire W19299;
wire W19300;
wire W19301;
wire W19302;
wire W19303;
wire W19304;
wire W19305;
wire W19306;
wire W19307;
wire W19308;
wire W19309;
wire W19310;
wire W19311;
wire W19312;
wire W19313;
wire W19314;
wire W19315;
wire W19316;
wire W19317;
wire W19318;
wire W19319;
wire W19320;
wire W19321;
wire W19322;
wire W19323;
wire W19324;
wire W19325;
wire W19326;
wire W19327;
wire W19328;
wire W19329;
wire W19330;
wire W19331;
wire W19332;
wire W19333;
wire W19334;
wire W19335;
wire W19336;
wire W19337;
wire W19338;
wire W19339;
wire W19340;
wire W19341;
wire W19342;
wire W19343;
wire W19344;
wire W19345;
wire W19346;
wire W19347;
wire W19348;
wire W19349;
wire W19350;
wire W19351;
wire W19352;
wire W19353;
wire W19354;
wire W19355;
wire W19356;
wire W19357;
wire W19358;
wire W19359;
wire W19360;
wire W19361;
wire W19362;
wire W19363;
wire W19364;
wire W19365;
wire W19366;
wire W19367;
wire W19368;
wire W19369;
wire W19370;
wire W19371;
wire W19372;
wire W19373;
wire W19374;
wire W19375;
wire W19376;
wire W19377;
wire W19378;
wire W19379;
wire W19380;
wire W19381;
wire W19382;
wire W19383;
wire W19384;
wire W19385;
wire W19386;
wire W19387;
wire W19388;
wire W19389;
wire W19390;
wire W19391;
wire W19392;
wire W19393;
wire W19394;
wire W19395;
wire W19396;
wire W19397;
wire W19398;
wire W19399;
wire W19400;
wire W19401;
wire W19402;
wire W19403;
wire W19404;
wire W19405;
wire W19406;
wire W19407;
wire W19408;
wire W19409;
wire W19410;
wire W19411;
wire W19412;
wire W19413;
wire W19414;
wire W19415;
wire W19416;
wire W19417;
wire W19418;
wire W19419;
wire W19420;
wire W19421;
wire W19422;
wire W19423;
wire W19424;
wire W19425;
wire W19426;
wire W19427;
wire W19428;
wire W19429;
wire W19430;
wire W19431;
wire W19432;
wire W19433;
wire W19434;
wire W19435;
wire W19436;
wire W19437;
wire W19438;
wire W19439;
wire W19440;
wire W19441;
wire W19442;
wire W19443;
wire W19444;
wire W19445;
wire W19446;
wire W19447;
wire W19448;
wire W19449;
wire W19450;
wire W19451;
wire W19452;
wire W19453;
wire W19454;
wire W19455;
wire W19456;
wire W19457;
wire W19458;
wire W19459;
wire W19460;
wire W19461;
wire W19462;
wire W19463;
wire W19464;
wire W19465;
wire W19466;
wire W19467;
wire W19468;
wire W19469;
wire W19470;
wire W19471;
wire W19472;
wire W19473;
wire W19474;
wire W19475;
wire W19476;
wire W19477;
wire W19478;
wire W19479;
wire W19480;
wire W19481;
wire W19482;
wire W19483;
wire W19484;
wire W19485;
wire W19486;
wire W19487;
wire W19488;
wire W19489;
wire W19490;
wire W19491;
wire W19492;
wire W19493;
wire W19494;
wire W19495;
wire W19496;
wire W19497;
wire W19498;
wire W19499;
wire W19500;
wire W19501;
wire W19502;
wire W19503;
wire W19504;
wire W19505;
wire W19506;
wire W19507;
wire W19508;
wire W19509;
wire W19510;
wire W19511;
wire W19512;
wire W19513;
wire W19514;
wire W19515;
wire W19516;
wire W19517;
wire W19518;
wire W19519;
wire W19520;
wire W19521;
wire W19522;
wire W19523;
wire W19524;
wire W19525;
wire W19526;
wire W19527;
wire W19528;
wire W19529;
wire W19530;
wire W19531;
wire W19532;
wire W19533;
wire W19534;
wire W19535;
wire W19536;
wire W19537;
wire W19538;
wire W19539;
wire W19540;
wire W19541;
wire W19542;
wire W19543;
wire W19544;
wire W19545;
wire W19546;
wire W19547;
wire W19548;
wire W19549;
wire W19550;
wire W19551;
wire W19552;
wire W19553;
wire W19554;
wire W19555;
wire W19556;
wire W19557;
wire W19558;
wire W19559;
wire W19560;
wire W19561;
wire W19562;
wire W19563;
wire W19564;
wire W19565;
wire W19566;
wire W19567;
wire W19568;
wire W19569;
wire W19570;
wire W19571;
wire W19572;
wire W19573;
wire W19574;
wire W19575;
wire W19576;
wire W19577;
wire W19578;
wire W19579;
wire W19580;
wire W19581;
wire W19582;
wire W19583;
wire W19584;
wire W19585;
wire W19586;
wire W19587;
wire W19588;
wire W19589;
wire W19590;
wire W19591;
wire W19592;
wire W19593;
wire W19594;
wire W19595;
wire W19596;
wire W19597;
wire W19598;
wire W19599;
wire W19600;
wire W19601;
wire W19602;
wire W19603;
wire W19604;
wire W19605;
wire W19606;
wire W19607;
wire W19608;
wire W19609;
wire W19610;
wire W19611;
wire W19612;
wire W19613;
wire W19614;
wire W19615;
wire W19616;
wire W19617;
wire W19618;
wire W19619;
wire W19620;
wire W19621;
wire W19622;
wire W19623;
wire W19624;
wire W19625;
wire W19626;
wire W19627;
wire W19628;
wire W19629;
wire W19630;
wire W19631;
wire W19632;
wire W19633;
wire W19634;
wire W19635;
wire W19636;
wire W19637;
wire W19638;
wire W19639;
wire W19640;
wire W19641;
wire W19642;
wire W19643;
wire W19644;
wire W19645;
wire W19646;
wire W19647;
wire W19648;
wire W19649;
wire W19650;
wire W19651;
wire W19652;
wire W19653;
wire W19654;
wire W19655;
wire W19656;
wire W19657;
wire W19658;
wire W19659;
wire W19660;
wire W19661;
wire W19662;
wire W19663;
wire W19664;
wire W19665;
wire W19666;
wire W19667;
wire W19668;
wire W19669;
wire W19670;
wire W19671;
wire W19672;
wire W19673;
wire W19674;
wire W19675;
wire W19676;
wire W19677;
wire W19678;
wire W19679;
wire W19680;
wire W19681;
wire W19682;
wire W19683;
wire W19684;
wire W19685;
wire W19686;
wire W19687;
wire W19688;
wire W19689;
wire W19690;
wire W19691;
wire W19692;
wire W19693;
wire W19694;
wire W19695;
wire W19696;
wire W19697;
wire W19698;
wire W19699;
wire W19700;
wire W19701;
wire W19702;
wire W19703;
wire W19704;
wire W19705;
wire W19706;
wire W19707;
wire W19708;
wire W19709;
wire W19710;
wire W19711;
wire W19712;
wire W19713;
wire W19714;
wire W19715;
wire W19716;
wire W19717;
wire W19718;
wire W19719;
wire W19720;
wire W19721;
wire W19722;
wire W19723;
wire W19724;
wire W19725;
wire W19726;
wire W19727;
wire W19728;
wire W19729;
wire W19730;
wire W19731;
wire W19732;
wire W19733;
wire W19734;
wire W19735;
wire W19736;
wire W19737;
wire W19738;
wire W19739;
wire W19740;
wire W19741;
wire W19742;
wire W19743;
wire W19744;
wire W19745;
wire W19746;
wire W19747;
wire W19748;
wire W19749;
wire W19750;
wire W19751;
wire W19752;
wire W19753;
wire W19754;
wire W19755;
wire W19756;
wire W19757;
wire W19758;
wire W19759;
wire W19760;
wire W19761;
wire W19762;
wire W19763;
wire W19764;
wire W19765;
wire W19766;
wire W19767;
wire W19768;
wire W19769;
wire W19770;
wire W19771;
wire W19772;
wire W19773;
wire W19774;
wire W19775;
wire W19776;
wire W19777;
wire W19778;
wire W19779;
wire W19780;
wire W19781;
wire W19782;
wire W19783;
wire W19784;
wire W19785;
wire W19786;
wire W19787;
wire W19788;
wire W19789;
wire W19790;
wire W19791;
wire W19792;
wire W19793;
wire W19794;
wire W19795;
wire W19796;
wire W19797;
wire W19798;
wire W19799;
wire W19800;
wire W19801;
wire W19802;
wire W19803;
wire W19804;
wire W19805;
wire W19806;
wire W19807;
wire W19808;
wire W19809;
wire W19810;
wire W19811;
wire W19812;
wire W19813;
wire W19814;
wire W19815;
wire W19816;
wire W19817;
wire W19818;
wire W19819;
wire W19820;
wire W19821;
wire W19822;
wire W19823;
wire W19824;
wire W19825;
wire W19826;
wire W19827;
wire W19828;
wire W19829;
wire W19830;
wire W19831;
wire W19832;
wire W19833;
wire W19834;
wire W19835;
wire W19836;
wire W19837;
wire W19838;
wire W19839;
wire W19840;
wire W19841;
wire W19842;
wire W19843;
wire W19844;
wire W19845;
wire W19846;
wire W19847;
wire W19848;
wire W19849;
wire W19850;
wire W19851;
wire W19852;
wire W19853;
wire W19854;
wire W19855;
wire W19856;
wire W19857;
wire W19858;
wire W19859;
wire W19860;
wire W19861;
wire W19862;
wire W19863;
wire W19864;
wire W19865;
wire W19866;
wire W19867;
wire W19868;
wire W19869;
wire W19870;
wire W19871;
wire W19872;
wire W19873;
wire W19874;
wire W19875;
wire W19876;
wire W19877;
wire W19878;
wire W19879;
wire W19880;
wire W19881;
wire W19882;
wire W19883;
wire W19884;
wire W19885;
wire W19886;
wire W19887;
wire W19888;
wire W19889;
wire W19890;
wire W19891;
wire W19892;
wire W19893;
wire W19894;
wire W19895;
wire W19896;
wire W19897;
wire W19898;
wire W19899;
wire W19900;
wire W19901;
wire W19902;
wire W19903;
wire W19904;
wire W19905;
wire W19906;
wire W19907;
wire W19908;
wire W19909;
wire W19910;
wire W19911;
wire W19912;
wire W19913;
wire W19914;
wire W19915;
wire W19916;
wire W19917;
wire W19918;
wire W19919;
wire W19920;
wire W19921;
wire W19922;
wire W19923;
wire W19924;
wire W19925;
wire W19926;
wire W19927;
wire W19928;
wire W19929;
wire W19930;
wire W19931;
wire W19932;
wire W19933;
wire W19934;
wire W19935;
wire W19936;
wire W19937;
wire W19938;
wire W19939;
wire W19940;
wire W19941;
wire W19942;
wire W19943;
wire W19944;
wire W19945;
wire W19946;
wire W19947;
wire W19948;
wire W19949;
wire W19950;
wire W19951;
wire W19952;
wire W19953;
wire W19954;
wire W19955;
wire W19956;
wire W19957;
wire W19958;
wire W19959;
wire W19960;
wire W19961;
wire W19962;
wire W19963;
wire W19964;
wire W19965;
wire W19966;
wire W19967;
wire W19968;
wire W19969;
wire W19970;
wire W19971;
wire W19972;
wire W19973;
wire W19974;
wire W19975;
wire W19976;
wire W19977;
wire W19978;
wire W19979;
wire W19980;
wire W19981;
wire W19982;
wire W19983;
wire W19984;
wire W19985;
wire W19986;
wire W19987;
wire W19988;
wire W19989;
wire W19990;
wire W19991;
wire W19992;
wire W19993;
wire W19994;
wire W19995;
wire W19996;
wire W19997;
wire W19998;
wire W19999;
wire W20000;
wire W20001;
wire W20002;
wire W20003;
wire W20004;
wire W20005;
wire W20006;
wire W20007;
wire W20008;
wire W20009;
wire W20010;
wire W20011;
wire W20012;
wire W20013;
wire W20014;
wire W20015;
wire W20016;
wire W20017;
wire W20018;
wire W20019;
wire W20020;
wire W20021;
wire W20022;
wire W20023;
wire W20024;
wire W20025;
wire W20026;
wire W20027;
wire W20028;
wire W20029;
wire W20030;
wire W20031;
wire W20032;
wire W20033;
wire W20034;
wire W20035;
wire W20036;
wire W20037;
wire W20038;
wire W20039;
wire W20040;
wire W20041;
wire W20042;
wire W20043;
wire W20044;
wire W20045;
wire W20046;
wire W20047;
wire W20048;
wire W20049;
wire W20050;
wire W20051;
wire W20052;
wire W20053;
wire W20054;
wire W20055;
wire W20056;
wire W20057;
wire W20058;
wire W20059;
wire W20060;
wire W20061;
wire W20062;
wire W20063;
wire W20064;
wire W20065;
wire W20066;
wire W20067;
wire W20068;
wire W20069;
wire W20070;
wire W20071;
wire W20072;
wire W20073;
wire W20074;
wire W20075;
wire W20076;
wire W20077;
wire W20078;
wire W20079;
wire W20080;
wire W20081;
wire W20082;
wire W20083;
wire W20084;
wire W20085;
wire W20086;
wire W20087;
wire W20088;
wire W20089;
wire W20090;
wire W20091;
wire W20092;
wire W20093;
wire W20094;
wire W20095;
wire W20096;
wire W20097;
wire W20098;
wire W20099;
wire W20100;
wire W20101;
wire W20102;
wire W20103;
wire W20104;
wire W20105;
wire W20106;
wire W20107;
wire W20108;
wire W20109;
wire W20110;
wire W20111;
wire W20112;
wire W20113;
wire W20114;
wire W20115;
wire W20116;
wire W20117;
wire W20118;
wire W20119;
wire W20120;
wire W20121;
wire W20122;
wire W20123;
wire W20124;
wire W20125;
wire W20126;
wire W20127;
wire W20128;
wire W20129;
wire W20130;
wire W20131;
wire W20132;
wire W20133;
wire W20134;
wire W20135;
wire W20136;
wire W20137;
wire W20138;
wire W20139;
wire W20140;
wire W20141;
wire W20142;
wire W20143;
wire W20144;
wire W20145;
wire W20146;
wire W20147;
wire W20148;
wire W20149;
wire W20150;
wire W20151;
wire W20152;
wire W20153;
wire W20154;
wire W20155;
wire W20156;
wire W20157;
wire W20158;
wire W20159;
wire W20160;
wire W20161;
wire W20162;
wire W20163;
wire W20164;
wire W20165;
wire W20166;
wire W20167;
wire W20168;
wire W20169;
wire W20170;
wire W20171;
wire W20172;
wire W20173;
wire W20174;
wire W20175;
wire W20176;
wire W20177;
wire W20178;
wire W20179;
wire W20180;
wire W20181;
wire W20182;
wire W20183;
wire W20184;
wire W20185;
wire W20186;
wire W20187;
wire W20188;
wire W20189;
wire W20190;
wire W20191;
wire W20192;
wire W20193;
wire W20194;
wire W20195;
wire W20196;
wire W20197;
wire W20198;
wire W20199;
wire W20200;
wire W20201;
wire W20202;
wire W20203;
wire W20204;
wire W20205;
wire W20206;
wire W20207;
wire W20208;
wire W20209;
wire W20210;
wire W20211;
wire W20212;
wire W20213;
wire W20214;
wire W20215;
wire W20216;
wire W20217;
wire W20218;
wire W20219;
wire W20220;
wire W20221;
wire W20222;
wire W20223;
wire W20224;
wire W20225;
wire W20226;
wire W20227;
wire W20228;
wire W20229;
wire W20230;
wire W20231;
wire W20232;
wire W20233;
wire W20234;
wire W20235;
wire W20236;
wire W20237;
wire W20238;
wire W20239;
wire W20240;
wire W20241;
wire W20242;
wire W20243;
wire W20244;
wire W20245;
wire W20246;
wire W20247;
wire W20248;
wire W20249;
wire W20250;
wire W20251;
wire W20252;
wire W20253;
wire W20254;
wire W20255;
wire W20256;
wire W20257;
wire W20258;
wire W20259;
wire W20260;
wire W20261;
wire W20262;
wire W20263;
wire W20264;
wire W20265;
wire W20266;
wire W20267;
wire W20268;
wire W20269;
wire W20270;
wire W20271;
wire W20272;
wire W20273;
wire W20274;
wire W20275;
wire W20276;
wire W20277;
wire W20278;
wire W20279;
wire W20280;
wire W20281;
wire W20282;
wire W20283;
wire W20284;
wire W20285;
wire W20286;
wire W20287;
wire W20288;
wire W20289;
wire W20290;
wire W20291;
wire W20292;
wire W20293;
wire W20294;
wire W20295;
wire W20296;
wire W20297;
wire W20298;
wire W20299;
wire W20300;
wire W20301;
wire W20302;
wire W20303;
wire W20304;
wire W20305;
wire W20306;
wire W20307;
wire W20308;
wire W20309;
wire W20310;
wire W20311;
wire W20312;
wire W20313;
wire W20314;
wire W20315;
wire W20316;
wire W20317;
wire W20318;
wire W20319;
wire W20320;
wire W20321;
wire W20322;
wire W20323;
wire W20324;
wire W20325;
wire W20326;
wire W20327;
wire W20328;
wire W20329;
wire W20330;

not G1 (O1, W1);
not G2 (O2, W2);
not G3 (O3, W3);
not G4 (O4, W4);
not G5 (O5, W5);
not G6 (O6, W6);
not G7 (O7, W7);
not G8 (O8, W8);
not G9 (O9, W9);
not G10 (O10, W10);
not G11 (O11, W11);
not G12 (O12, W12);
not G13 (O13, W13);
not G14 (O14, W14);
not G15 (O15, W15);
not G16 (O16, W16);
not G17 (O17, W17);
not G18 (O18, W18);
not G19 (O19, W19);
not G20 (O20, W20);
not G21 (O21, W21);
not G22 (O22, W22);
not G23 (O23, W23);
not G24 (O24, W24);
not G25 (O25, W25);
not G26 (O26, W26);
not G27 (O27, W27);
not G28 (O28, W28);
not G29 (O29, W29);
not G30 (O30, W30);
not G31 (O31, W31);
not G32 (O32, W32);
not G33 (O33, W33);
not G34 (O34, W34);
not G35 (O35, W35);
not G36 (O36, W36);
not G37 (O37, W37);
not G38 (O38, W38);
not G39 (O39, W39);
not G40 (O40, W40);
not G41 (O41, W41);
not G42 (O42, W42);
not G43 (O43, W43);
not G44 (O44, W44);
not G45 (O45, W45);
not G46 (O46, W46);
not G47 (O47, W47);
not G48 (O48, W48);
not G49 (O49, W49);
not G50 (O50, W50);
not G51 (O51, W51);
not G52 (O52, W52);
not G53 (O53, W53);
not G54 (O54, W54);
not G55 (O55, W55);
not G56 (O56, W56);
not G57 (O57, W57);
not G58 (O58, W58);
not G59 (O59, W59);
not G60 (O60, W60);
not G61 (O61, W61);
not G62 (O62, W62);
not G63 (O63, W63);
not G64 (O64, W64);
not G65 (O65, W65);
not G66 (O66, W66);
not G67 (O67, W67);
not G68 (O68, W68);
not G69 (O69, W69);
not G70 (O70, W70);
not G71 (O71, W71);
not G72 (O72, W72);
not G73 (O73, W73);
not G74 (O74, W74);
not G75 (O75, W75);
not G76 (O76, W76);
not G77 (O77, W77);
not G78 (O78, W78);
not G79 (O79, W79);
not G80 (O80, W80);
not G81 (O81, W81);
not G82 (O82, W82);
not G83 (O83, W83);
not G84 (O84, W84);
not G85 (O85, W85);
not G86 (O86, W86);
not G87 (O87, W87);
not G88 (O88, W88);
not G89 (O89, W89);
not G90 (O90, W90);
not G91 (O91, W91);
not G92 (O92, W92);
not G93 (O93, W93);
not G94 (O94, W94);
not G95 (O95, W95);
not G96 (O96, W96);
not G97 (O97, W97);
not G98 (O98, W98);
not G99 (O99, W99);
not G100 (O100, W100);
not G101 (O101, W101);
not G102 (O102, W102);
not G103 (O103, W103);
not G104 (O104, W104);
not G105 (O105, W105);
not G106 (O106, W106);
not G107 (O107, W107);
not G108 (O108, W108);
not G109 (O109, W109);
not G110 (O110, W110);
not G111 (O111, W111);
not G112 (O112, W112);
not G113 (O113, W113);
not G114 (O114, W114);
not G115 (O115, W115);
not G116 (O116, W116);
not G117 (O117, W117);
not G118 (O118, W118);
not G119 (O119, W119);
not G120 (O120, W120);
not G121 (O121, W121);
not G122 (O122, W122);
not G123 (O123, W123);
not G124 (O124, W124);
not G125 (O125, W125);
not G126 (O126, W126);
not G127 (O127, W127);
not G128 (O128, W128);
not G129 (O129, W129);
not G130 (O130, W130);
not G131 (O131, W131);
not G132 (O132, W132);
not G133 (O133, W133);
not G134 (O134, W134);
not G135 (O135, W135);
not G136 (O136, W136);
not G137 (O137, W137);
not G138 (O138, W138);
not G139 (O139, W139);
not G140 (O140, W140);
not G141 (O141, W141);
not G142 (O142, W142);
not G143 (O143, W143);
not G144 (O144, W144);
not G145 (O145, W145);
not G146 (O146, W146);
not G147 (O147, W147);
not G148 (O148, W148);
not G149 (O149, W149);
not G150 (O150, W150);
not G151 (O151, W151);
not G152 (O152, W152);
not G153 (O153, W153);
not G154 (O154, W154);
not G155 (O155, W155);
not G156 (O156, W156);
not G157 (O157, W157);
not G158 (O158, W158);
not G159 (O159, W159);
not G160 (O160, W160);
not G161 (O161, W161);
not G162 (O162, W162);
not G163 (O163, W163);
not G164 (O164, W164);
not G165 (O165, W165);
not G166 (O166, W166);
not G167 (O167, W167);
not G168 (O168, W168);
not G169 (O169, W169);
not G170 (O170, W170);
not G171 (O171, W171);
not G172 (O172, W172);
not G173 (O173, W173);
not G174 (O174, W174);
not G175 (O175, W175);
not G176 (O176, W176);
not G177 (O177, W177);
not G178 (O178, W178);
not G179 (O179, W179);
not G180 (O180, W180);
not G181 (O181, W181);
not G182 (O182, W182);
not G183 (O183, W183);
not G184 (O184, W184);
not G185 (O185, W185);
not G186 (O186, W186);
not G187 (O187, W187);
not G188 (O188, W188);
not G189 (O189, W189);
not G190 (O190, W190);
not G191 (O191, W191);
not G192 (O192, W192);
not G193 (O193, W193);
not G194 (O194, W194);
not G195 (O195, W195);
not G196 (O196, W196);
not G197 (O197, W197);
not G198 (O198, W198);
not G199 (O199, W199);
not G200 (O200, W200);
not G201 (O201, W201);
not G202 (O202, W202);
not G203 (O203, W203);
not G204 (O204, W204);
not G205 (O205, W205);
not G206 (O206, W206);
not G207 (O207, W207);
not G208 (O208, W208);
not G209 (O209, W209);
not G210 (O210, W210);
not G211 (O211, W211);
not G212 (O212, W212);
not G213 (O213, W213);
not G214 (O214, W214);
not G215 (O215, W215);
not G216 (O216, W216);
not G217 (O217, W217);
not G218 (O218, W218);
not G219 (O219, W219);
not G220 (O220, W220);
not G221 (O221, W221);
not G222 (O222, W222);
not G223 (O223, W223);
not G224 (O224, W224);
not G225 (O225, W225);
not G226 (O226, W226);
not G227 (O227, W227);
not G228 (O228, W228);
not G229 (O229, W229);
not G230 (O230, W230);
not G231 (O231, W231);
not G232 (O232, W232);
not G233 (O233, W233);
not G234 (O234, W234);
not G235 (O235, W235);
not G236 (O236, W236);
not G237 (O237, W237);
not G238 (O238, W238);
not G239 (O239, W239);
not G240 (O240, W240);
not G241 (O241, W241);
not G242 (O242, W242);
not G243 (O243, W243);
not G244 (O244, W244);
not G245 (O245, W245);
not G246 (O246, W246);
not G247 (O247, W247);
not G248 (O248, W248);
not G249 (O249, W249);
not G250 (O250, W250);
not G251 (O251, W251);
not G252 (O252, W252);
not G253 (O253, W253);
not G254 (O254, W254);
not G255 (O255, W255);
not G256 (O256, W256);
not G257 (O257, W257);
not G258 (O258, W258);
not G259 (O259, W259);
not G260 (O260, W260);
not G261 (O261, W261);
not G262 (O262, W262);
not G263 (O263, W263);
not G264 (O264, W264);
not G265 (O265, W265);
not G266 (O266, W266);
not G267 (O267, W267);
not G268 (O268, W268);
not G269 (O269, W269);
not G270 (O270, W270);
not G271 (O271, W271);
not G272 (O272, W272);
not G273 (O273, W273);
not G274 (O274, W274);
not G275 (O275, W275);
not G276 (O276, W276);
not G277 (O277, W277);
not G278 (O278, W278);
not G279 (O279, W279);
not G280 (O280, W280);
not G281 (O281, W281);
not G282 (O282, W282);
not G283 (O283, W283);
not G284 (O284, W284);
not G285 (O285, W285);
not G286 (O286, W286);
not G287 (O287, W287);
not G288 (O288, W288);
not G289 (O289, W289);
not G290 (O290, W290);
not G291 (O291, W291);
not G292 (O292, W292);
not G293 (O293, W293);
not G294 (O294, W294);
not G295 (O295, W295);
not G296 (O296, W296);
not G297 (O297, W297);
not G298 (O298, W298);
not G299 (O299, W299);
not G300 (O300, W300);
not G301 (O301, W301);
not G302 (O302, W302);
not G303 (O303, W303);
not G304 (O304, W304);
not G305 (O305, W305);
not G306 (O306, W306);
not G307 (O307, W307);
not G308 (O308, W308);
not G309 (O309, W309);
not G310 (O310, W310);
not G311 (O311, W311);
not G312 (O312, W312);
not G313 (O313, W313);
not G314 (O314, W314);
not G315 (O315, W315);
not G316 (O316, W316);
not G317 (O317, W317);
not G318 (O318, W318);
not G319 (O319, W319);
not G320 (O320, W320);
not G321 (O321, W321);
not G322 (O322, W322);
not G323 (O323, W323);
not G324 (O324, W324);
not G325 (O325, W325);
not G326 (O326, W326);
not G327 (O327, W327);
not G328 (O328, W328);
not G329 (O329, W329);
not G330 (O330, W330);
not G331 (O331, W331);
not G332 (O332, W332);
not G333 (O333, W333);
not G334 (O334, W334);
not G335 (O335, W335);
not G336 (O336, W336);
not G337 (O337, W337);
not G338 (O338, W338);
not G339 (O339, W339);
not G340 (O340, W340);
not G341 (O341, W341);
not G342 (O342, W342);
not G343 (O343, W343);
not G344 (O344, W344);
not G345 (O345, W345);
not G346 (O346, W346);
not G347 (O347, W347);
not G348 (O348, W348);
not G349 (O349, W349);
not G350 (O350, W350);
not G351 (O351, W351);
not G352 (O352, W352);
not G353 (O353, W353);
not G354 (O354, W354);
not G355 (O355, W355);
not G356 (O356, W356);
not G357 (O357, W357);
not G358 (O358, W358);
not G359 (O359, W359);
not G360 (O360, W360);
not G361 (O361, W361);
not G362 (O362, W362);
not G363 (O363, W363);
not G364 (O364, W364);
not G365 (O365, W365);
not G366 (O366, W366);
not G367 (O367, W367);
not G368 (O368, W368);
not G369 (O369, W369);
not G370 (O370, W370);
not G371 (O371, W371);
not G372 (O372, W372);
not G373 (O373, W373);
not G374 (O374, W374);
not G375 (O375, W375);
not G376 (O376, W376);
not G377 (O377, W377);
not G378 (O378, W378);
not G379 (O379, W379);
not G380 (O380, W380);
not G381 (O381, W381);
not G382 (O382, W382);
not G383 (O383, W383);
not G384 (O384, W384);
not G385 (O385, W385);
not G386 (O386, W386);
not G387 (O387, W387);
not G388 (O388, W388);
not G389 (O389, W389);
not G390 (O390, W390);
not G391 (O391, W391);
not G392 (O392, W392);
not G393 (O393, W393);
not G394 (O394, W394);
not G395 (O395, W395);
not G396 (O396, W396);
not G397 (O397, W397);
not G398 (O398, W398);
not G399 (O399, W399);
not G400 (O400, W400);
not G401 (O401, W401);
not G402 (O402, W402);
not G403 (O403, W403);
not G404 (O404, W404);
not G405 (O405, W405);
not G406 (O406, W406);
not G407 (O407, W407);
not G408 (O408, W408);
not G409 (O409, W409);
not G410 (O410, W410);
not G411 (O411, W411);
not G412 (O412, W412);
not G413 (O413, W413);
not G414 (O414, W414);
not G415 (O415, W415);
not G416 (O416, W416);
not G417 (O417, W417);
not G418 (O418, W418);
not G419 (O419, W419);
not G420 (O420, W420);
not G421 (O421, W421);
not G422 (O422, W422);
not G423 (O423, W423);
not G424 (O424, W424);
not G425 (O425, W425);
not G426 (O426, W426);
not G427 (O427, W427);
not G428 (O428, W428);
not G429 (O429, W429);
not G430 (O430, W430);
not G431 (O431, W431);
not G432 (O432, W432);
not G433 (O433, W433);
not G434 (O434, W434);
not G435 (O435, W435);
not G436 (O436, W436);
not G437 (O437, W437);
not G438 (O438, W438);
not G439 (O439, W439);
not G440 (O440, W440);
not G441 (O441, W441);
not G442 (O442, W442);
not G443 (O443, W443);
not G444 (O444, W444);
not G445 (O445, W445);
not G446 (O446, W446);
not G447 (O447, W447);
not G448 (O448, W448);
not G449 (O449, W449);
not G450 (O450, W450);
not G451 (O451, W451);
not G452 (O452, W452);
not G453 (O453, W453);
not G454 (O454, W454);
not G455 (O455, W455);
not G456 (O456, W456);
not G457 (O457, W457);
not G458 (O458, W458);
not G459 (O459, W459);
not G460 (O460, W460);
not G461 (O461, W461);
not G462 (O462, W462);
not G463 (O463, W463);
not G464 (O464, W464);
not G465 (O465, W465);
not G466 (O466, W466);
not G467 (O467, W467);
not G468 (O468, W468);
not G469 (O469, W469);
not G470 (O470, W470);
not G471 (O471, W471);
not G472 (O472, W472);
not G473 (O473, W473);
not G474 (O474, W474);
not G475 (O475, W475);
not G476 (O476, W476);
not G477 (O477, W477);
not G478 (O478, W478);
not G479 (O479, W479);
not G480 (O480, W480);
not G481 (O481, W481);
not G482 (O482, W482);
not G483 (O483, W483);
not G484 (O484, W484);
not G485 (O485, W485);
not G486 (O486, W486);
not G487 (O487, W487);
not G488 (O488, W488);
not G489 (O489, W489);
not G490 (O490, W490);
not G491 (O491, W491);
not G492 (O492, W492);
not G493 (O493, W493);
not G494 (O494, W494);
not G495 (O495, W495);
not G496 (O496, W496);
not G497 (O497, W497);
not G498 (O498, W498);
not G499 (O499, W499);
not G500 (O500, W500);
not G501 (O501, W501);
not G502 (O502, W502);
not G503 (O503, W503);
not G504 (O504, W504);
not G505 (O505, W505);
not G506 (O506, W506);
not G507 (O507, W507);
not G508 (O508, W508);
not G509 (O509, W509);
not G510 (O510, W510);
not G511 (O511, W511);
not G512 (O512, W512);
not G513 (O513, W513);
not G514 (O514, W514);
not G515 (O515, W515);
not G516 (O516, W516);
not G517 (O517, W517);
not G518 (O518, W518);
not G519 (O519, W519);
not G520 (O520, W520);
not G521 (O521, W521);
not G522 (O522, W522);
not G523 (O523, W523);
not G524 (O524, W524);
not G525 (O525, W525);
not G526 (O526, W526);
not G527 (O527, W527);
not G528 (O528, W528);
not G529 (O529, W529);
not G530 (O530, W530);
not G531 (O531, W531);
not G532 (O532, W532);
not G533 (O533, W533);
not G534 (O534, W534);
not G535 (O535, W535);
not G536 (O536, W536);
not G537 (O537, W537);
not G538 (O538, W538);
not G539 (O539, W539);
not G540 (O540, W540);
not G541 (O541, W541);
not G542 (O542, W542);
not G543 (O543, W543);
not G544 (O544, W544);
not G545 (O545, W545);
not G546 (O546, W546);
not G547 (O547, W547);
not G548 (O548, W548);
not G549 (O549, W549);
not G550 (O550, W550);
not G551 (O551, W551);
not G552 (O552, W552);
not G553 (O553, W553);
not G554 (O554, W554);
not G555 (O555, W555);
not G556 (O556, W556);
not G557 (O557, W557);
not G558 (O558, W558);
not G559 (O559, W559);
not G560 (O560, W560);
not G561 (O561, W561);
not G562 (O562, W562);
not G563 (O563, W563);
not G564 (O564, W564);
not G565 (O565, W565);
not G566 (O566, W566);
not G567 (O567, W567);
not G568 (O568, W568);
not G569 (O569, W569);
not G570 (O570, W570);
not G571 (O571, W571);
not G572 (O572, W572);
not G573 (O573, W573);
not G574 (O574, W574);
not G575 (O575, W575);
not G576 (O576, W576);
not G577 (O577, W577);
not G578 (O578, W578);
not G579 (O579, W579);
not G580 (O580, W580);
not G581 (O581, W581);
not G582 (O582, W582);
not G583 (O583, W583);
not G584 (O584, W584);
not G585 (O585, W585);
not G586 (O586, W586);
not G587 (O587, W587);
not G588 (O588, W588);
not G589 (O589, W589);
not G590 (O590, W590);
not G591 (O591, W591);
not G592 (O592, W592);
not G593 (O593, W593);
not G594 (O594, W594);
not G595 (O595, W595);
not G596 (O596, W596);
not G597 (O597, W597);
not G598 (O598, W598);
not G599 (O599, W599);
not G600 (O600, W600);
not G601 (O601, W601);
not G602 (O602, W602);
not G603 (O603, W603);
not G604 (O604, W604);
not G605 (O605, W605);
not G606 (O606, W606);
not G607 (O607, W607);
not G608 (O608, W608);
not G609 (O609, W609);
not G610 (O610, W610);
not G611 (O611, W611);
not G612 (O612, W612);
not G613 (O613, W613);
not G614 (O614, W614);
not G615 (O615, W615);
not G616 (O616, W616);
not G617 (O617, W617);
not G618 (O618, W618);
not G619 (O619, W619);
not G620 (O620, W620);
not G621 (O621, W621);
not G622 (O622, W622);
not G623 (O623, W623);
not G624 (O624, W624);
not G625 (O625, W625);
not G626 (O626, W626);
not G627 (O627, W627);
not G628 (O628, W628);
not G629 (O629, W629);
not G630 (O630, W630);
not G631 (O631, W631);
not G632 (O632, W632);
not G633 (O633, W633);
not G634 (O634, W634);
not G635 (O635, W635);
not G636 (O636, W636);
not G637 (O637, W637);
not G638 (O638, W638);
not G639 (O639, W639);
not G640 (O640, W640);
not G641 (O641, W641);
not G642 (O642, W642);
not G643 (O643, W643);
not G644 (O644, W644);
not G645 (O645, W645);
not G646 (O646, W646);
not G647 (O647, W647);
not G648 (O648, W648);
not G649 (O649, W649);
not G650 (O650, W650);
not G651 (O651, W651);
not G652 (O652, W652);
not G653 (O653, W653);
not G654 (O654, W654);
not G655 (O655, W655);
not G656 (O656, W656);
not G657 (O657, W657);
not G658 (O658, W658);
not G659 (O659, W659);
not G660 (O660, W660);
not G661 (O661, W661);
not G662 (O662, W662);
not G663 (O663, W663);
not G664 (O664, W664);
not G665 (O665, W665);
not G666 (O666, W666);
not G667 (O667, W667);
not G668 (O668, W668);
not G669 (O669, W669);
not G670 (O670, W670);
not G671 (O671, W671);
not G672 (O672, W672);
not G673 (O673, W673);
not G674 (O674, W674);
not G675 (O675, W675);
not G676 (O676, W676);
not G677 (O677, W677);
not G678 (O678, W678);
not G679 (O679, W679);
not G680 (O680, W680);
not G681 (O681, W681);
not G682 (O682, W682);
not G683 (O683, W683);
not G684 (O684, W684);
not G685 (O685, W685);
not G686 (O686, W686);
not G687 (O687, W687);
not G688 (O688, W688);
not G689 (O689, W689);
not G690 (O690, W690);
not G691 (O691, W691);
not G692 (O692, W692);
not G693 (O693, W693);
not G694 (O694, W694);
not G695 (O695, W695);
not G696 (O696, W696);
not G697 (O697, W697);
not G698 (O698, W698);
not G699 (O699, W699);
not G700 (O700, W700);
not G701 (O701, W701);
not G702 (O702, W702);
not G703 (O703, W703);
not G704 (O704, W704);
not G705 (O705, W705);
not G706 (O706, W706);
not G707 (O707, W707);
not G708 (O708, W708);
not G709 (O709, W709);
not G710 (O710, W710);
not G711 (O711, W711);
not G712 (O712, W712);
not G713 (O713, W713);
not G714 (O714, W714);
not G715 (O715, W715);
not G716 (O716, W716);
not G717 (O717, W717);
not G718 (O718, W718);
not G719 (O719, W719);
not G720 (O720, W720);
not G721 (O721, W721);
not G722 (O722, W722);
not G723 (O723, W723);
not G724 (O724, W724);
not G725 (O725, W725);
not G726 (O726, W726);
not G727 (O727, W727);
not G728 (O728, W728);
not G729 (O729, W729);
not G730 (O730, W730);
not G731 (O731, W731);
not G732 (O732, W732);
not G733 (O733, W733);
not G734 (O734, W734);
not G735 (O735, W735);
not G736 (O736, W736);
not G737 (O737, W737);
not G738 (O738, W738);
not G739 (O739, W739);
not G740 (O740, W740);
not G741 (O741, W741);
not G742 (O742, W742);
not G743 (O743, W743);
not G744 (O744, W744);
not G745 (O745, W745);
not G746 (O746, W746);
not G747 (O747, W747);
not G748 (O748, W748);
not G749 (O749, W749);
not G750 (O750, W750);
not G751 (O751, W751);
not G752 (O752, W752);
not G753 (O753, W753);
not G754 (O754, W754);
not G755 (O755, W755);
not G756 (O756, W756);
not G757 (O757, W757);
not G758 (O758, W758);
not G759 (O759, W759);
not G760 (O760, W760);
not G761 (O761, W761);
not G762 (O762, W762);
not G763 (O763, W763);
not G764 (O764, W764);
not G765 (O765, W765);
not G766 (O766, W766);
not G767 (O767, W767);
not G768 (O768, W768);
not G769 (O769, W769);
not G770 (O770, W770);
not G771 (O771, W771);
not G772 (O772, W772);
not G773 (O773, W773);
not G774 (O774, W774);
not G775 (O775, W775);
not G776 (O776, W776);
not G777 (O777, W777);
not G778 (O778, W778);
not G779 (O779, W779);
not G780 (O780, W780);
not G781 (O781, W781);
not G782 (O782, W782);
not G783 (O783, W783);
not G784 (O784, W784);
not G785 (O785, W785);
not G786 (O786, W786);
not G787 (O787, W787);
not G788 (O788, W788);
not G789 (O789, W789);
not G790 (O790, W790);
not G791 (O791, W791);
not G792 (O792, W792);
not G793 (O793, W793);
not G794 (O794, W794);
not G795 (O795, W795);
not G796 (O796, W796);
not G797 (O797, W797);
not G798 (O798, W798);
not G799 (O799, W799);
not G800 (O800, W800);
not G801 (O801, W801);
not G802 (O802, W802);
not G803 (O803, W803);
not G804 (O804, W804);
not G805 (O805, W805);
not G806 (O806, W806);
not G807 (O807, W807);
not G808 (O808, W808);
not G809 (O809, W809);
not G810 (O810, W810);
not G811 (O811, W811);
not G812 (O812, W812);
not G813 (O813, W813);
not G814 (O814, W814);
not G815 (O815, W815);
not G816 (O816, W816);
not G817 (O817, W817);
not G818 (O818, W818);
not G819 (O819, W819);
not G820 (O820, W820);
not G821 (O821, W821);
not G822 (O822, W822);
not G823 (O823, W823);
not G824 (O824, W824);
not G825 (O825, W825);
not G826 (O826, W826);
not G827 (O827, W827);
not G828 (O828, W828);
not G829 (O829, W829);
not G830 (O830, W830);
not G831 (O831, W831);
not G832 (O832, W832);
not G833 (O833, W833);
not G834 (O834, W834);
not G835 (O835, W835);
not G836 (O836, W836);
not G837 (O837, W837);
not G838 (O838, W838);
not G839 (O839, W839);
not G840 (O840, W840);
not G841 (O841, W841);
not G842 (O842, W842);
not G843 (O843, W843);
not G844 (O844, W844);
not G845 (O845, W845);
not G846 (O846, W846);
not G847 (O847, W847);
not G848 (O848, W848);
not G849 (O849, W849);
not G850 (O850, W850);
not G851 (O851, W851);
not G852 (O852, W852);
not G853 (O853, W853);
not G854 (O854, W854);
not G855 (O855, W855);
not G856 (O856, W856);
not G857 (O857, W857);
not G858 (O858, W858);
not G859 (O859, W859);
not G860 (O860, W860);
not G861 (O861, W861);
not G862 (O862, W862);
not G863 (O863, W863);
not G864 (O864, W864);
not G865 (O865, W865);
not G866 (O866, W866);
not G867 (O867, W867);
not G868 (O868, W868);
not G869 (O869, W869);
not G870 (O870, W870);
not G871 (O871, W871);
not G872 (O872, W872);
not G873 (O873, W873);
not G874 (O874, W874);
not G875 (O875, W875);
not G876 (O876, W876);
not G877 (O877, W877);
not G878 (O878, W878);
not G879 (O879, W879);
not G880 (O880, W880);
not G881 (O881, W881);
not G882 (O882, W882);
not G883 (O883, W883);
not G884 (O884, W884);
not G885 (O885, W885);
not G886 (O886, W886);
not G887 (O887, W887);
not G888 (O888, W888);
not G889 (O889, W889);
not G890 (O890, W890);
not G891 (O891, W891);
not G892 (O892, W892);
not G893 (O893, W893);
not G894 (O894, W894);
not G895 (O895, W895);
not G896 (O896, W896);
not G897 (O897, W897);
not G898 (O898, W898);
not G899 (O899, W899);
not G900 (O900, W900);
not G901 (O901, W901);
not G902 (O902, W902);
not G903 (O903, W903);
not G904 (O904, W904);
not G905 (O905, W905);
not G906 (O906, W906);
not G907 (O907, W907);
not G908 (O908, W908);
not G909 (O909, W909);
not G910 (O910, W910);
not G911 (O911, W911);
not G912 (O912, W912);
not G913 (O913, W913);
not G914 (O914, W914);
not G915 (O915, W915);
not G916 (O916, W916);
not G917 (O917, W917);
not G918 (O918, W918);
not G919 (O919, W919);
not G920 (O920, W920);
not G921 (O921, W921);
not G922 (O922, W922);
not G923 (O923, W923);
not G924 (O924, W924);
not G925 (O925, W925);
not G926 (O926, W926);
not G927 (O927, W927);
not G928 (O928, W928);
not G929 (O929, W929);
not G930 (O930, W930);
not G931 (O931, W931);
not G932 (O932, W932);
not G933 (O933, W933);
not G934 (O934, W934);
not G935 (O935, W935);
not G936 (O936, W936);
not G937 (O937, W937);
not G938 (O938, W938);
not G939 (O939, W939);
not G940 (O940, W940);
not G941 (O941, W941);
not G942 (O942, W942);
not G943 (O943, W943);
not G944 (O944, W944);
not G945 (O945, W945);
not G946 (O946, W946);
not G947 (O947, W947);
not G948 (O948, W948);
not G949 (O949, W949);
not G950 (O950, W950);
not G951 (O951, W951);
not G952 (O952, W952);
not G953 (O953, W953);
not G954 (O954, W954);
not G955 (O955, W955);
not G956 (O956, W956);
not G957 (O957, W957);
not G958 (O958, W958);
not G959 (O959, W959);
not G960 (O960, W960);
not G961 (O961, W961);
not G962 (O962, W962);
not G963 (O963, W963);
not G964 (O964, W964);
not G965 (O965, W965);
not G966 (O966, W966);
not G967 (O967, W967);
not G968 (O968, W968);
not G969 (O969, W969);
not G970 (O970, W970);
not G971 (O971, W971);
not G972 (O972, W972);
not G973 (O973, W973);
not G974 (O974, W974);
not G975 (O975, W975);
not G976 (O976, W976);
not G977 (O977, W977);
not G978 (O978, W978);
not G979 (O979, W979);
not G980 (O980, W980);
not G981 (O981, W981);
not G982 (O982, W982);
not G983 (O983, W983);
not G984 (O984, W984);
not G985 (O985, W985);
not G986 (O986, W986);
not G987 (O987, W987);
not G988 (O988, W988);
not G989 (O989, W989);
not G990 (O990, W990);
not G991 (O991, W991);
not G992 (O992, W992);
not G993 (O993, W993);
not G994 (O994, W994);
not G995 (O995, W995);
not G996 (O996, W996);
not G997 (O997, W997);
not G998 (O998, W998);
not G999 (O999, W999);
not G1000 (O1000, W1000);
not G1001 (O1001, W1001);
not G1002 (O1002, W1002);
not G1003 (O1003, W1003);
not G1004 (O1004, W1004);
not G1005 (O1005, W1005);
not G1006 (O1006, W1006);
not G1007 (O1007, W1007);
not G1008 (O1008, W1008);
not G1009 (O1009, W1009);
not G1010 (O1010, W1010);
not G1011 (O1011, W1011);
not G1012 (O1012, W1012);
not G1013 (O1013, W1013);
not G1014 (O1014, W1014);
not G1015 (O1015, W1015);
not G1016 (O1016, W1016);
not G1017 (O1017, W1017);
not G1018 (O1018, W1018);
not G1019 (O1019, W1019);
not G1020 (O1020, W1020);
not G1021 (O1021, W1021);
not G1022 (O1022, W1022);
not G1023 (O1023, W1023);
not G1024 (O1024, W1024);
not G1025 (O1025, W1025);
not G1026 (O1026, W1026);
not G1027 (O1027, W1027);
not G1028 (O1028, W1028);
not G1029 (O1029, W1029);
not G1030 (O1030, W1030);
not G1031 (O1031, W1031);
not G1032 (O1032, W1032);
not G1033 (O1033, W1033);
not G1034 (O1034, W1034);
not G1035 (O1035, W1035);
not G1036 (O1036, W1036);
not G1037 (O1037, W1037);
not G1038 (O1038, W1038);
not G1039 (O1039, W1039);
not G1040 (O1040, W1040);
not G1041 (O1041, W1041);
not G1042 (O1042, W1042);
not G1043 (O1043, W1043);
not G1044 (O1044, W1044);
not G1045 (O1045, W1045);
not G1046 (O1046, W1046);
not G1047 (O1047, W1047);
not G1048 (O1048, W1048);
not G1049 (O1049, W1049);
not G1050 (O1050, W1050);
not G1051 (O1051, W1051);
not G1052 (O1052, W1052);
not G1053 (O1053, W1053);
not G1054 (O1054, W1054);
not G1055 (O1055, W1055);
not G1056 (O1056, W1056);
not G1057 (O1057, W1057);
not G1058 (O1058, W1058);
not G1059 (O1059, W1059);
not G1060 (O1060, W1060);
not G1061 (O1061, W1061);
not G1062 (O1062, W1062);
not G1063 (O1063, W1063);
not G1064 (O1064, W1064);
not G1065 (O1065, W1065);
not G1066 (O1066, W1066);
not G1067 (O1067, W1067);
not G1068 (O1068, W1068);
not G1069 (O1069, W1069);
not G1070 (O1070, W1070);
not G1071 (O1071, W1071);
not G1072 (O1072, W1072);
not G1073 (O1073, W1073);
not G1074 (O1074, W1074);
not G1075 (O1075, W1075);
not G1076 (O1076, W1076);
not G1077 (O1077, W1077);
not G1078 (O1078, W1078);
not G1079 (O1079, W1079);
not G1080 (O1080, W1080);
not G1081 (O1081, W1081);
not G1082 (O1082, W1082);
not G1083 (O1083, W1083);
not G1084 (O1084, W1084);
not G1085 (O1085, W1085);
not G1086 (O1086, W1086);
not G1087 (O1087, W1087);
not G1088 (O1088, W1088);
not G1089 (O1089, W1089);
not G1090 (O1090, W1090);
not G1091 (O1091, W1091);
not G1092 (O1092, W1092);
not G1093 (O1093, W1093);
not G1094 (O1094, W1094);
not G1095 (O1095, W1095);
not G1096 (O1096, W1096);
not G1097 (O1097, W1097);
not G1098 (O1098, W1098);
not G1099 (O1099, W1099);
not G1100 (O1100, W1100);
not G1101 (O1101, W1101);
not G1102 (O1102, W1102);
not G1103 (O1103, W1103);
not G1104 (O1104, W1104);
not G1105 (O1105, W1105);
not G1106 (O1106, W1106);
not G1107 (O1107, W1107);
not G1108 (O1108, W1108);
not G1109 (O1109, W1109);
not G1110 (O1110, W1110);
not G1111 (O1111, W1111);
not G1112 (O1112, W1112);
not G1113 (O1113, W1113);
not G1114 (O1114, W1114);
not G1115 (O1115, W1115);
not G1116 (O1116, W1116);
not G1117 (O1117, W1117);
not G1118 (O1118, W1118);
not G1119 (O1119, W1119);
not G1120 (O1120, W1120);
not G1121 (O1121, W1121);
not G1122 (O1122, W1122);
not G1123 (O1123, W1123);
not G1124 (O1124, W1124);
not G1125 (O1125, W1125);
not G1126 (O1126, W1126);
not G1127 (O1127, W1127);
not G1128 (O1128, W1128);
not G1129 (O1129, W1129);
not G1130 (O1130, W1130);
not G1131 (O1131, W1131);
not G1132 (O1132, W1132);
not G1133 (O1133, W1133);
not G1134 (O1134, W1134);
not G1135 (O1135, W1135);
not G1136 (O1136, W1136);
not G1137 (O1137, W1137);
not G1138 (O1138, W1138);
not G1139 (O1139, W1139);
not G1140 (O1140, W1140);
not G1141 (O1141, W1141);
not G1142 (O1142, W1142);
not G1143 (O1143, W1143);
not G1144 (O1144, W1144);
not G1145 (O1145, W1145);
not G1146 (O1146, W1146);
not G1147 (O1147, W1147);
not G1148 (O1148, W1148);
not G1149 (O1149, W1149);
not G1150 (O1150, W1150);
not G1151 (O1151, W1151);
not G1152 (O1152, W1152);
not G1153 (O1153, W1153);
not G1154 (O1154, W1154);
not G1155 (O1155, W1155);
not G1156 (O1156, W1156);
not G1157 (O1157, W1157);
not G1158 (O1158, W1158);
not G1159 (O1159, W1159);
not G1160 (O1160, W1160);
not G1161 (O1161, W1161);
not G1162 (O1162, W1162);
not G1163 (O1163, W1163);
not G1164 (O1164, W1164);
not G1165 (O1165, W1165);
not G1166 (O1166, W1166);
not G1167 (O1167, W1167);
not G1168 (O1168, W1168);
not G1169 (O1169, W1169);
not G1170 (O1170, W1170);
not G1171 (O1171, W1171);
not G1172 (O1172, W1172);
not G1173 (O1173, W1173);
not G1174 (O1174, W1174);
not G1175 (O1175, W1175);
not G1176 (O1176, W1176);
not G1177 (O1177, W1177);
not G1178 (O1178, W1178);
not G1179 (O1179, W1179);
not G1180 (O1180, W1180);
not G1181 (O1181, W1181);
not G1182 (O1182, W1182);
not G1183 (O1183, W1183);
not G1184 (O1184, W1184);
not G1185 (O1185, W1185);
not G1186 (O1186, W1186);
not G1187 (O1187, W1187);
not G1188 (O1188, W1188);
not G1189 (O1189, W1189);
not G1190 (O1190, W1190);
not G1191 (O1191, W1191);
not G1192 (O1192, W1192);
not G1193 (O1193, W1193);
not G1194 (O1194, W1194);
not G1195 (O1195, W1195);
not G1196 (O1196, W1196);
not G1197 (O1197, W1197);
not G1198 (O1198, W1198);
not G1199 (O1199, W1199);
not G1200 (O1200, W1200);
not G1201 (O1201, W1201);
not G1202 (O1202, W1202);
not G1203 (O1203, W1203);
not G1204 (O1204, W1204);
not G1205 (O1205, W1205);
not G1206 (O1206, W1206);
not G1207 (O1207, W1207);
not G1208 (O1208, W1208);
not G1209 (O1209, W1209);
not G1210 (O1210, W1210);
not G1211 (O1211, W1211);
not G1212 (O1212, W1212);
not G1213 (O1213, W1213);
not G1214 (O1214, W1214);
not G1215 (O1215, W1215);
not G1216 (O1216, W1216);
not G1217 (O1217, W1217);
not G1218 (O1218, W1218);
not G1219 (O1219, W1219);
not G1220 (O1220, W1220);
not G1221 (O1221, W1221);
not G1222 (O1222, W1222);
not G1223 (O1223, W1223);
not G1224 (O1224, W1224);
not G1225 (O1225, W1225);
not G1226 (O1226, W1226);
not G1227 (O1227, W1227);
not G1228 (O1228, W1228);
not G1229 (O1229, W1229);
not G1230 (O1230, W1230);
not G1231 (O1231, W1231);
not G1232 (O1232, W1232);
not G1233 (O1233, W1233);
not G1234 (O1234, W1234);
not G1235 (O1235, W1235);
not G1236 (O1236, W1236);
not G1237 (O1237, W1237);
not G1238 (O1238, W1238);
not G1239 (O1239, W1239);
not G1240 (O1240, W1240);
not G1241 (O1241, W1241);
not G1242 (O1242, W1242);
not G1243 (O1243, W1243);
not G1244 (O1244, W1244);
not G1245 (O1245, W1245);
not G1246 (O1246, W1246);
not G1247 (O1247, W1247);
not G1248 (O1248, W1248);
not G1249 (O1249, W1249);
not G1250 (O1250, W1250);
not G1251 (O1251, W1251);
not G1252 (O1252, W1252);
not G1253 (O1253, W1253);
not G1254 (O1254, W1254);
not G1255 (O1255, W1255);
not G1256 (O1256, W1256);
not G1257 (O1257, W1257);
not G1258 (O1258, W1258);
not G1259 (O1259, W1259);
not G1260 (O1260, W1260);
not G1261 (O1261, W1261);
not G1262 (O1262, W1262);
not G1263 (O1263, W1263);
not G1264 (O1264, W1264);
not G1265 (O1265, W1265);
not G1266 (O1266, W1266);
not G1267 (O1267, W1267);
not G1268 (O1268, W1268);
not G1269 (O1269, W1269);
not G1270 (O1270, W1270);
not G1271 (O1271, W1271);
not G1272 (O1272, W1272);
not G1273 (O1273, W1273);
not G1274 (O1274, W1274);
not G1275 (O1275, W1275);
not G1276 (O1276, W1276);
not G1277 (O1277, W1277);
not G1278 (O1278, W1278);
not G1279 (O1279, W1279);
not G1280 (O1280, W1280);
not G1281 (O1281, W1281);
not G1282 (O1282, W1282);
not G1283 (O1283, W1283);
not G1284 (O1284, W1284);
not G1285 (O1285, W1285);
not G1286 (O1286, W1286);
not G1287 (O1287, W1287);
not G1288 (O1288, W1288);
not G1289 (O1289, W1289);
not G1290 (O1290, W1290);
not G1291 (O1291, W1291);
not G1292 (O1292, W1292);
not G1293 (O1293, W1293);
not G1294 (O1294, W1294);
not G1295 (O1295, W1295);
not G1296 (O1296, W1296);
not G1297 (O1297, W1297);
not G1298 (O1298, W1298);
not G1299 (O1299, W1299);
not G1300 (O1300, W1300);
not G1301 (O1301, W1301);
not G1302 (O1302, W1302);
not G1303 (O1303, W1303);
not G1304 (O1304, W1304);
not G1305 (O1305, W1305);
not G1306 (O1306, W1306);
not G1307 (O1307, W1307);
not G1308 (O1308, W1308);
not G1309 (O1309, W1309);
not G1310 (O1310, W1310);
not G1311 (O1311, W1311);
not G1312 (O1312, W1312);
not G1313 (O1313, W1313);
not G1314 (O1314, W1314);
not G1315 (O1315, W1315);
not G1316 (O1316, W1316);
not G1317 (O1317, W1317);
not G1318 (O1318, W1318);
not G1319 (O1319, W1319);
not G1320 (O1320, W1320);
not G1321 (O1321, W1321);
not G1322 (O1322, W1322);
not G1323 (O1323, W1323);
not G1324 (O1324, W1324);
not G1325 (O1325, W1325);
not G1326 (O1326, W1326);
not G1327 (O1327, W1327);
not G1328 (O1328, W1328);
not G1329 (O1329, W1329);
not G1330 (O1330, W1330);
not G1331 (O1331, W1331);
not G1332 (O1332, W1332);
not G1333 (O1333, W1333);
not G1334 (O1334, W1334);
not G1335 (O1335, W1335);
not G1336 (O1336, W1336);
not G1337 (O1337, W1337);
not G1338 (O1338, W1338);
not G1339 (O1339, W1339);
not G1340 (O1340, W1340);
not G1341 (O1341, W1341);
not G1342 (O1342, W1342);
not G1343 (O1343, W1343);
not G1344 (O1344, W1344);
not G1345 (O1345, W1345);
not G1346 (O1346, W1346);
not G1347 (O1347, W1347);
not G1348 (O1348, W1348);
not G1349 (O1349, W1349);
not G1350 (O1350, W1350);
not G1351 (O1351, W1351);
not G1352 (O1352, W1352);
not G1353 (O1353, W1353);
not G1354 (O1354, W1354);
not G1355 (O1355, W1355);
not G1356 (O1356, W1356);
not G1357 (O1357, W1357);
not G1358 (O1358, W1358);
not G1359 (O1359, W1359);
not G1360 (O1360, W1360);
not G1361 (O1361, W1361);
not G1362 (O1362, W1362);
not G1363 (O1363, W1363);
not G1364 (O1364, W1364);
not G1365 (O1365, W1365);
not G1366 (O1366, W1366);
not G1367 (O1367, W1367);
not G1368 (O1368, W1368);
not G1369 (O1369, W1369);
not G1370 (O1370, W1370);
not G1371 (O1371, W1371);
not G1372 (O1372, W1372);
not G1373 (O1373, W1373);
not G1374 (O1374, W1374);
not G1375 (O1375, W1375);
not G1376 (O1376, W1376);
not G1377 (O1377, W1377);
not G1378 (O1378, W1378);
not G1379 (O1379, W1379);
not G1380 (O1380, W1380);
not G1381 (O1381, W1381);
not G1382 (O1382, W1382);
not G1383 (O1383, W1383);
not G1384 (O1384, W1384);
not G1385 (O1385, W1385);
not G1386 (O1386, W1386);
not G1387 (O1387, W1387);
not G1388 (O1388, W1388);
not G1389 (O1389, W1389);
not G1390 (O1390, W1390);
not G1391 (O1391, W1391);
not G1392 (O1392, W1392);
not G1393 (O1393, W1393);
not G1394 (O1394, W1394);
not G1395 (O1395, W1395);
not G1396 (O1396, W1396);
not G1397 (O1397, W1397);
not G1398 (W1, W1398);
not G1399 (W2, W1399);
not G1400 (W3, W1400);
not G1401 (W4, W1401);
not G1402 (W5, W1402);
not G1403 (W6, W1403);
not G1404 (W7, W1404);
not G1405 (W8, W1405);
not G1406 (W9, W1406);
not G1407 (W10, W1407);
not G1408 (W11, W1408);
not G1409 (W12, W1409);
not G1410 (W13, W1410);
not G1411 (W14, W1411);
not G1412 (W15, W1412);
not G1413 (W16, W1413);
not G1414 (W17, W1414);
not G1415 (W18, W1415);
not G1416 (W19, W1416);
not G1417 (W20, W1417);
not G1418 (W21, W1418);
not G1419 (W22, W1419);
not G1420 (W23, W1420);
not G1421 (W24, W1421);
not G1422 (W25, W1422);
not G1423 (W26, W1423);
not G1424 (W27, W1424);
not G1425 (W28, W1425);
not G1426 (W29, W1426);
not G1427 (W30, W1427);
not G1428 (W31, W1428);
not G1429 (W32, W1429);
not G1430 (W33, W1430);
not G1431 (W34, W1431);
not G1432 (W35, W1432);
not G1433 (W36, W1433);
not G1434 (W37, W1434);
not G1435 (W38, W1435);
not G1436 (W39, W1436);
not G1437 (W40, W1437);
not G1438 (W41, W1438);
not G1439 (W42, W1439);
not G1440 (W43, W1440);
not G1441 (W44, W1441);
not G1442 (W45, W1442);
not G1443 (W46, W1443);
not G1444 (W47, W1444);
not G1445 (W48, W1445);
not G1446 (W49, W1446);
not G1447 (W50, W1447);
not G1448 (W51, W1448);
not G1449 (W52, W1449);
not G1450 (W53, W1450);
not G1451 (W54, W1451);
not G1452 (W55, W1452);
not G1453 (W56, W1453);
not G1454 (W57, W1454);
not G1455 (W58, W1455);
not G1456 (W59, W1456);
not G1457 (W60, W1457);
not G1458 (W61, W1458);
not G1459 (W62, W1459);
not G1460 (W63, W1460);
not G1461 (W64, W1461);
not G1462 (W65, W1462);
not G1463 (W66, W1463);
not G1464 (W67, W1464);
not G1465 (W68, W1465);
not G1466 (W69, W1466);
not G1467 (W70, W1467);
not G1468 (W71, W1468);
not G1469 (W72, W1469);
not G1470 (W73, W1470);
not G1471 (W74, W1471);
not G1472 (W75, W1472);
not G1473 (W76, W1473);
not G1474 (W77, W1474);
not G1475 (W78, W1475);
not G1476 (W79, W1476);
not G1477 (W80, W1477);
not G1478 (W81, W1478);
not G1479 (W82, W1479);
not G1480 (W83, W1480);
not G1481 (W84, W1481);
not G1482 (W85, W1482);
not G1483 (W86, W1483);
not G1484 (W87, W1484);
not G1485 (W88, W1485);
not G1486 (W89, W1486);
not G1487 (W90, W1487);
not G1488 (W91, W1488);
not G1489 (W92, W1489);
not G1490 (W93, W1490);
not G1491 (W94, W1491);
not G1492 (W95, W1492);
not G1493 (W96, W1493);
not G1494 (W97, W1494);
not G1495 (W98, W1495);
not G1496 (W99, W1496);
not G1497 (W100, W1497);
not G1498 (W101, W1498);
not G1499 (W102, W1499);
not G1500 (W103, W1500);
not G1501 (W104, W1501);
not G1502 (W105, W1502);
not G1503 (W106, W1503);
not G1504 (W107, W1504);
not G1505 (W108, W1505);
not G1506 (W109, W1506);
not G1507 (W110, W1507);
not G1508 (W111, W1508);
not G1509 (W112, W1509);
not G1510 (W113, W1510);
not G1511 (W114, W1511);
not G1512 (W115, W1512);
not G1513 (W116, W1513);
not G1514 (W117, W1514);
not G1515 (W118, W1515);
not G1516 (W119, W1516);
not G1517 (W120, W1517);
not G1518 (W121, W1518);
not G1519 (W122, W1519);
not G1520 (W123, W1520);
not G1521 (W124, W1521);
not G1522 (W125, W1522);
not G1523 (W126, W1523);
not G1524 (W127, W1524);
not G1525 (W128, W1525);
not G1526 (W129, W1526);
not G1527 (W130, W1527);
not G1528 (W131, W1528);
not G1529 (W132, W1529);
not G1530 (W133, W1530);
not G1531 (W134, W1531);
not G1532 (W135, W1532);
not G1533 (W136, W1533);
not G1534 (W137, W1534);
not G1535 (W138, W1535);
not G1536 (W139, W1536);
not G1537 (W140, W1537);
not G1538 (W141, W1538);
not G1539 (W142, W1539);
not G1540 (W143, W1540);
not G1541 (W144, W1541);
not G1542 (W145, W1542);
not G1543 (W146, W1543);
not G1544 (W147, W1544);
not G1545 (W148, W1545);
not G1546 (W149, W1546);
not G1547 (W150, W1547);
not G1548 (W151, W1548);
not G1549 (W152, W1549);
not G1550 (W153, W1550);
not G1551 (W154, W1551);
not G1552 (W155, W1552);
not G1553 (W156, W1553);
not G1554 (W157, W1554);
not G1555 (W158, W1555);
not G1556 (W159, W1556);
not G1557 (W160, W1557);
not G1558 (W161, W1558);
not G1559 (W162, W1559);
not G1560 (W163, W1560);
not G1561 (W164, W1561);
not G1562 (W165, W1562);
not G1563 (W166, W1563);
not G1564 (W167, W1564);
not G1565 (W168, W1565);
not G1566 (W169, W1566);
not G1567 (W170, W1567);
not G1568 (W171, W1568);
not G1569 (W172, W1569);
not G1570 (W173, W1570);
not G1571 (W174, W1571);
not G1572 (W175, W1572);
not G1573 (W176, W1573);
not G1574 (W177, W1574);
not G1575 (W178, W1575);
not G1576 (W179, W1576);
not G1577 (W180, W1577);
not G1578 (W181, W1578);
not G1579 (W182, W1579);
not G1580 (W183, W1580);
not G1581 (W184, W1581);
not G1582 (W185, W1582);
not G1583 (W186, W1583);
not G1584 (W187, W1584);
not G1585 (W188, W1585);
not G1586 (W189, W1586);
not G1587 (W190, W1587);
not G1588 (W191, W1588);
not G1589 (W192, W1589);
not G1590 (W193, W1590);
not G1591 (W194, W1591);
not G1592 (W195, W1592);
not G1593 (W196, W1593);
not G1594 (W197, W1594);
not G1595 (W198, W1595);
not G1596 (W199, W1596);
not G1597 (W200, W1597);
not G1598 (W201, W1598);
not G1599 (W202, W1599);
not G1600 (W203, W1600);
not G1601 (W204, W1601);
not G1602 (W205, W1602);
not G1603 (W206, W1603);
not G1604 (W207, W1604);
not G1605 (W208, W1605);
not G1606 (W209, W1606);
not G1607 (W210, W1607);
not G1608 (W211, W1608);
not G1609 (W212, W1609);
not G1610 (W213, W1610);
not G1611 (W214, W1611);
not G1612 (W215, W1612);
not G1613 (W216, W1613);
not G1614 (W217, W1614);
not G1615 (W218, W1615);
not G1616 (W219, W1616);
not G1617 (W220, W1617);
not G1618 (W221, W1618);
not G1619 (W222, W1619);
not G1620 (W223, W1620);
not G1621 (W224, W1621);
not G1622 (W225, W1622);
not G1623 (W226, W1623);
not G1624 (W227, W1624);
not G1625 (W228, W1625);
not G1626 (W229, W1626);
not G1627 (W230, W1627);
not G1628 (W231, W1628);
not G1629 (W232, W1629);
not G1630 (W233, W1630);
not G1631 (W234, W1631);
not G1632 (W235, W1632);
not G1633 (W236, W1633);
not G1634 (W237, W1634);
not G1635 (W238, W1635);
not G1636 (W239, W1636);
not G1637 (W240, W1637);
not G1638 (W241, W1638);
not G1639 (W242, W1639);
not G1640 (W243, W1640);
not G1641 (W244, W1641);
not G1642 (W245, W1642);
not G1643 (W246, W1643);
not G1644 (W247, W1644);
not G1645 (W248, W1645);
not G1646 (W249, W1646);
not G1647 (W250, W1647);
not G1648 (W251, W1648);
not G1649 (W252, W1649);
not G1650 (W253, W1650);
not G1651 (W254, W1651);
not G1652 (W255, W1652);
not G1653 (W256, W1653);
not G1654 (W257, W1654);
not G1655 (W258, W1655);
not G1656 (W259, W1656);
not G1657 (W260, W1657);
not G1658 (W261, W1658);
not G1659 (W262, W1659);
not G1660 (W263, W1660);
not G1661 (W264, W1661);
not G1662 (W265, W1662);
not G1663 (W266, W1663);
not G1664 (W267, W1664);
not G1665 (W268, W1665);
not G1666 (W269, W1666);
not G1667 (W270, W1667);
not G1668 (W271, W1668);
not G1669 (W272, W1669);
not G1670 (W273, W1670);
not G1671 (W274, W1671);
not G1672 (W275, W1672);
not G1673 (W276, W1673);
not G1674 (W277, W1674);
not G1675 (W278, W1675);
not G1676 (W279, W1676);
not G1677 (W280, W1677);
not G1678 (W281, W1678);
not G1679 (W282, W1679);
not G1680 (W283, W1680);
not G1681 (W284, W1681);
not G1682 (W285, W1682);
not G1683 (W286, W1683);
not G1684 (W287, W1684);
not G1685 (W288, W1685);
not G1686 (W289, W1686);
not G1687 (W290, W1687);
not G1688 (W291, W1688);
not G1689 (W292, W1689);
not G1690 (W293, W1690);
not G1691 (W294, W1691);
not G1692 (W295, W1692);
not G1693 (W296, W1693);
not G1694 (W297, W1694);
not G1695 (W298, W1695);
not G1696 (W299, W1696);
not G1697 (W300, W1697);
not G1698 (W301, W1698);
not G1699 (W302, W1699);
not G1700 (W303, W1700);
not G1701 (W304, W1701);
not G1702 (W305, W1702);
not G1703 (W306, W1703);
not G1704 (W307, W1704);
not G1705 (W308, W1705);
not G1706 (W309, W1706);
not G1707 (W310, W1707);
not G1708 (W311, W1708);
not G1709 (W312, W1709);
not G1710 (W313, W1710);
not G1711 (W314, W1711);
not G1712 (W315, W1712);
not G1713 (W316, W1713);
not G1714 (W317, W1714);
not G1715 (W318, W1715);
not G1716 (W319, W1716);
not G1717 (W320, W1717);
not G1718 (W321, W1718);
not G1719 (W322, W1719);
not G1720 (W323, W1720);
not G1721 (W324, W1721);
not G1722 (W325, W1722);
not G1723 (W326, W1723);
not G1724 (W327, W1724);
not G1725 (W328, W1725);
not G1726 (W329, W1726);
not G1727 (W330, W1727);
not G1728 (W331, W1728);
not G1729 (W332, W1729);
not G1730 (W333, W1730);
not G1731 (W334, W1731);
not G1732 (W335, W1732);
not G1733 (W336, W1733);
not G1734 (W337, W1734);
not G1735 (W338, W1735);
not G1736 (W339, W1736);
not G1737 (W340, W1737);
not G1738 (W341, W1738);
not G1739 (W342, W1739);
not G1740 (W343, W1740);
not G1741 (W344, W1741);
not G1742 (W345, W1742);
not G1743 (W346, W1743);
not G1744 (W347, W1744);
not G1745 (W348, W1745);
not G1746 (W349, W1746);
not G1747 (W350, W1747);
not G1748 (W351, W1748);
not G1749 (W352, W1749);
not G1750 (W353, W1750);
not G1751 (W354, W1751);
not G1752 (W355, W1752);
not G1753 (W356, W1753);
not G1754 (W357, W1754);
not G1755 (W358, W1755);
not G1756 (W359, W1756);
not G1757 (W360, W1757);
not G1758 (W361, W1758);
not G1759 (W362, W1759);
not G1760 (W363, W1760);
not G1761 (W364, W1761);
not G1762 (W365, W1762);
not G1763 (W366, W1763);
not G1764 (W367, W1764);
not G1765 (W368, W1765);
not G1766 (W369, W1766);
not G1767 (W370, W1767);
not G1768 (W371, W1768);
not G1769 (W372, W1769);
not G1770 (W373, W1770);
not G1771 (W374, W1771);
not G1772 (W375, W1772);
not G1773 (W376, W1773);
not G1774 (W377, W1774);
not G1775 (W378, W1775);
not G1776 (W379, W1776);
not G1777 (W380, W1777);
not G1778 (W381, W1778);
not G1779 (W382, W1779);
not G1780 (W383, W1780);
not G1781 (W384, W1781);
not G1782 (W385, W1782);
not G1783 (W386, W1783);
not G1784 (W387, W1784);
not G1785 (W388, W1785);
not G1786 (W389, W1786);
not G1787 (W390, W1787);
not G1788 (W391, W1788);
not G1789 (W392, W1789);
not G1790 (W393, W1790);
not G1791 (W394, W1791);
not G1792 (W395, W1792);
not G1793 (W396, W1793);
not G1794 (W397, W1794);
not G1795 (W398, W1795);
not G1796 (W399, W1796);
not G1797 (W400, W1797);
not G1798 (W401, W1798);
not G1799 (W402, W1799);
not G1800 (W403, W1800);
not G1801 (W404, W1801);
not G1802 (W405, W1802);
not G1803 (W406, W1803);
not G1804 (W407, W1804);
not G1805 (W408, W1805);
not G1806 (W409, W1806);
not G1807 (W410, W1807);
not G1808 (W411, W1808);
not G1809 (W412, W1809);
not G1810 (W413, W1810);
not G1811 (W414, W1811);
not G1812 (W415, W1812);
not G1813 (W416, W1813);
not G1814 (W417, W1814);
not G1815 (W418, W1815);
not G1816 (W419, W1816);
not G1817 (W420, W1817);
not G1818 (W421, W1818);
not G1819 (W422, W1819);
not G1820 (W423, W1820);
not G1821 (W424, W1821);
not G1822 (W425, W1822);
not G1823 (W426, W1823);
not G1824 (W427, W1824);
not G1825 (W428, W1825);
not G1826 (W429, W1826);
not G1827 (W430, W1827);
not G1828 (W431, W1828);
not G1829 (W432, W1829);
not G1830 (W433, W1830);
not G1831 (W434, W1831);
not G1832 (W435, W1832);
not G1833 (W436, W1833);
not G1834 (W437, W1834);
not G1835 (W438, W1835);
not G1836 (W439, W1836);
not G1837 (W440, W1837);
not G1838 (W441, W1838);
not G1839 (W442, W1839);
not G1840 (W443, W1840);
not G1841 (W444, W1841);
not G1842 (W445, W1842);
not G1843 (W446, W1843);
not G1844 (W447, W1844);
not G1845 (W448, W1845);
not G1846 (W449, W1846);
not G1847 (W450, W1847);
not G1848 (W451, W1848);
not G1849 (W452, W1849);
not G1850 (W453, W1850);
not G1851 (W454, W1851);
not G1852 (W455, W1852);
not G1853 (W456, W1853);
not G1854 (W457, W1854);
not G1855 (W458, W1855);
not G1856 (W459, W1856);
not G1857 (W460, W1857);
not G1858 (W461, W1858);
not G1859 (W462, W1859);
not G1860 (W463, W1860);
not G1861 (W464, W1861);
not G1862 (W465, W1862);
not G1863 (W466, W1863);
not G1864 (W467, W1864);
not G1865 (W468, W1865);
not G1866 (W469, W1866);
not G1867 (W470, W1867);
not G1868 (W471, W1868);
not G1869 (W472, W1869);
not G1870 (W473, W1870);
not G1871 (W474, W1871);
not G1872 (W475, W1872);
not G1873 (W476, W1873);
not G1874 (W477, W1874);
not G1875 (W478, W1875);
not G1876 (W479, W1876);
not G1877 (W480, W1877);
not G1878 (W481, W1878);
not G1879 (W482, W1879);
not G1880 (W483, W1880);
not G1881 (W484, W1881);
not G1882 (W485, W1882);
not G1883 (W486, W1883);
not G1884 (W487, W1884);
not G1885 (W488, W1885);
not G1886 (W489, W1886);
not G1887 (W490, W1887);
not G1888 (W491, W1888);
not G1889 (W492, W1889);
not G1890 (W493, W1890);
not G1891 (W494, W1891);
not G1892 (W495, W1892);
not G1893 (W496, W1893);
not G1894 (W497, W1894);
not G1895 (W498, W1895);
not G1896 (W499, W1896);
not G1897 (W500, W1897);
not G1898 (W501, W1898);
not G1899 (W502, W1899);
not G1900 (W503, W1900);
not G1901 (W504, W1901);
not G1902 (W505, W1902);
not G1903 (W506, W1903);
not G1904 (W507, W1904);
not G1905 (W508, W1905);
not G1906 (W509, W1906);
not G1907 (W510, W1907);
not G1908 (W511, W1908);
not G1909 (W512, W1909);
not G1910 (W513, W1910);
not G1911 (W514, W1911);
not G1912 (W515, W1912);
not G1913 (W516, W1913);
not G1914 (W517, W1914);
not G1915 (W518, W1915);
not G1916 (W519, W1916);
not G1917 (W520, W1917);
not G1918 (W521, W1918);
not G1919 (W522, W1919);
not G1920 (W523, W1920);
not G1921 (W524, W1921);
not G1922 (W525, W1922);
not G1923 (W526, W1923);
not G1924 (W527, W1924);
not G1925 (W528, W1925);
not G1926 (W529, W1926);
not G1927 (W530, W1927);
not G1928 (W531, W1928);
not G1929 (W532, W1929);
not G1930 (W533, W1930);
not G1931 (W534, W1931);
not G1932 (W535, W1932);
not G1933 (W536, W1933);
not G1934 (W537, W1934);
not G1935 (W538, W1935);
not G1936 (W539, W1936);
not G1937 (W540, W1937);
not G1938 (W541, W1938);
not G1939 (W542, W1939);
not G1940 (W543, W1940);
not G1941 (W544, W1941);
not G1942 (W545, W1942);
not G1943 (W546, W1943);
not G1944 (W547, W1944);
not G1945 (W548, W1945);
not G1946 (W549, W1946);
not G1947 (W550, W1947);
not G1948 (W551, W1948);
not G1949 (W552, W1949);
not G1950 (W553, W1950);
not G1951 (W554, W1951);
not G1952 (W555, W1952);
not G1953 (W556, W1953);
not G1954 (W557, W1954);
not G1955 (W558, W1955);
not G1956 (W559, W1956);
not G1957 (W560, W1957);
not G1958 (W561, W1958);
not G1959 (W562, W1959);
not G1960 (W563, W1960);
not G1961 (W564, W1961);
not G1962 (W565, W1962);
not G1963 (W566, W1963);
not G1964 (W567, W1964);
not G1965 (W568, W1965);
not G1966 (W569, W1966);
not G1967 (W570, W1967);
not G1968 (W571, W1968);
not G1969 (W572, W1969);
not G1970 (W573, W1970);
not G1971 (W574, W1971);
not G1972 (W575, W1972);
not G1973 (W576, W1973);
not G1974 (W577, W1974);
not G1975 (W578, W1975);
not G1976 (W579, W1976);
not G1977 (W580, W1977);
not G1978 (W581, W1978);
not G1979 (W582, W1979);
not G1980 (W583, W1980);
not G1981 (W584, W1981);
not G1982 (W585, W1982);
not G1983 (W586, W1983);
not G1984 (W587, W1984);
not G1985 (W588, W1985);
not G1986 (W589, W1986);
not G1987 (W590, W1987);
not G1988 (W591, W1988);
not G1989 (W592, W1989);
not G1990 (W593, W1990);
not G1991 (W594, W1991);
not G1992 (W595, W1992);
not G1993 (W596, W1993);
not G1994 (W597, W1994);
not G1995 (W598, W1995);
not G1996 (W599, W1996);
not G1997 (W600, W1997);
not G1998 (W601, W1998);
not G1999 (W602, W1999);
not G2000 (W603, W2000);
not G2001 (W604, W2001);
not G2002 (W605, W2002);
not G2003 (W606, W2003);
not G2004 (W607, W2004);
not G2005 (W608, W2005);
not G2006 (W609, W2006);
not G2007 (W610, W2007);
not G2008 (W611, W2008);
not G2009 (W612, W2009);
not G2010 (W613, W2010);
not G2011 (W614, W2011);
not G2012 (W615, W2012);
not G2013 (W616, W2013);
not G2014 (W617, W2014);
not G2015 (W618, W2015);
not G2016 (W619, W2016);
not G2017 (W620, W2017);
not G2018 (W621, W2018);
not G2019 (W622, W2019);
not G2020 (W623, W2020);
not G2021 (W624, W2021);
not G2022 (W625, W2022);
not G2023 (W626, W2023);
not G2024 (W627, W2024);
not G2025 (W628, W2025);
not G2026 (W629, W2026);
not G2027 (W630, W2027);
not G2028 (W631, W2028);
not G2029 (W632, W2029);
not G2030 (W633, W2030);
not G2031 (W634, W2031);
not G2032 (W635, W2032);
not G2033 (W636, W2033);
not G2034 (W637, W2034);
not G2035 (W638, W2035);
not G2036 (W639, W2036);
not G2037 (W640, W2037);
not G2038 (W641, W2038);
not G2039 (W642, W2039);
not G2040 (W643, W2040);
not G2041 (W644, W2041);
not G2042 (W645, W2042);
not G2043 (W646, W2043);
not G2044 (W647, W2044);
not G2045 (W648, W2045);
not G2046 (W649, W2046);
not G2047 (W650, W2047);
not G2048 (W651, W2048);
not G2049 (W652, W2049);
not G2050 (W653, W2050);
not G2051 (W654, W2051);
not G2052 (W655, W2052);
not G2053 (W656, W2053);
not G2054 (W657, W2054);
not G2055 (W658, W2055);
not G2056 (W659, W2056);
not G2057 (W660, W2057);
not G2058 (W661, W2058);
not G2059 (W662, W2059);
not G2060 (W663, W2060);
not G2061 (W664, W2061);
not G2062 (W665, W2062);
not G2063 (W666, W2063);
not G2064 (W667, W2064);
not G2065 (W668, W2065);
not G2066 (W669, W2066);
not G2067 (W670, W2067);
not G2068 (W671, W2068);
not G2069 (W672, W2069);
not G2070 (W673, W2070);
not G2071 (W674, W2071);
not G2072 (W675, W2072);
not G2073 (W676, W2073);
not G2074 (W677, W2074);
not G2075 (W678, W2075);
not G2076 (W679, W2076);
not G2077 (W680, W2077);
not G2078 (W681, W2078);
not G2079 (W682, W2079);
not G2080 (W683, W2080);
not G2081 (W684, W2081);
not G2082 (W685, W2082);
not G2083 (W686, W2083);
not G2084 (W687, W2084);
not G2085 (W688, W2085);
not G2086 (W689, W2086);
not G2087 (W690, W2087);
not G2088 (W691, W2088);
not G2089 (W692, W2089);
not G2090 (W693, W2090);
not G2091 (W694, W2091);
not G2092 (W695, W2092);
not G2093 (W696, W2093);
not G2094 (W697, W2094);
not G2095 (W698, W2095);
not G2096 (W699, W2096);
not G2097 (W700, W2097);
not G2098 (W701, W2098);
not G2099 (W702, W2099);
not G2100 (W703, W2100);
not G2101 (W704, W2101);
not G2102 (W705, W2102);
not G2103 (W706, W2103);
not G2104 (W707, W2104);
not G2105 (W708, W2105);
not G2106 (W709, W2106);
not G2107 (W710, W2107);
not G2108 (W711, W2108);
not G2109 (W712, W2109);
not G2110 (W713, W2110);
not G2111 (W714, W2111);
not G2112 (W715, W2112);
not G2113 (W716, W2113);
not G2114 (W717, W2114);
not G2115 (W718, W2115);
not G2116 (W719, W2116);
not G2117 (W720, W2117);
not G2118 (W721, W2118);
not G2119 (W722, W2119);
not G2120 (W723, W2120);
not G2121 (W724, W2121);
not G2122 (W725, W2122);
not G2123 (W726, W2123);
not G2124 (W727, W2124);
not G2125 (W728, W2125);
not G2126 (W729, W2126);
not G2127 (W730, W2127);
not G2128 (W731, W2128);
not G2129 (W732, W2129);
not G2130 (W733, W2130);
not G2131 (W734, W2131);
not G2132 (W735, W2132);
not G2133 (W736, W2133);
not G2134 (W737, W2134);
not G2135 (W738, W2135);
not G2136 (W739, W2136);
not G2137 (W740, W2137);
not G2138 (W741, W2138);
not G2139 (W742, W2139);
not G2140 (W743, W2140);
not G2141 (W744, W2141);
not G2142 (W745, W2142);
not G2143 (W746, W2143);
not G2144 (W747, W2144);
not G2145 (W748, W2145);
not G2146 (W749, W2146);
not G2147 (W750, W2147);
not G2148 (W751, W2148);
not G2149 (W752, W2149);
not G2150 (W753, W2150);
not G2151 (W754, W2151);
not G2152 (W755, W2152);
not G2153 (W756, W2153);
not G2154 (W757, W2154);
not G2155 (W758, W2155);
not G2156 (W759, W2156);
not G2157 (W760, W2157);
not G2158 (W761, W2158);
not G2159 (W762, W2159);
not G2160 (W763, W2160);
not G2161 (W764, W2161);
not G2162 (W765, W2162);
not G2163 (W766, W2163);
not G2164 (W767, W2164);
not G2165 (W768, W2165);
not G2166 (W769, W2166);
not G2167 (W770, W2167);
not G2168 (W771, W2168);
not G2169 (W772, W2169);
not G2170 (W773, W2170);
not G2171 (W774, W2171);
not G2172 (W775, W2172);
not G2173 (W776, W2173);
not G2174 (W777, W2174);
not G2175 (W778, W2175);
not G2176 (W779, W2176);
not G2177 (W780, W2177);
not G2178 (W781, W2178);
not G2179 (W782, W2179);
not G2180 (W783, W2180);
not G2181 (W784, W2181);
not G2182 (W785, W2182);
not G2183 (W786, W2183);
not G2184 (W787, W2184);
not G2185 (W788, W2185);
not G2186 (W789, W2186);
not G2187 (W790, W2187);
not G2188 (W791, W2188);
not G2189 (W792, W2189);
not G2190 (W793, W2190);
not G2191 (W794, W2191);
not G2192 (W795, W2192);
not G2193 (W796, W2193);
not G2194 (W797, W2194);
not G2195 (W798, W2195);
not G2196 (W799, W2196);
not G2197 (W800, W2197);
not G2198 (W801, W2198);
not G2199 (W802, W2199);
not G2200 (W803, W2200);
not G2201 (W804, W2201);
not G2202 (W805, W2202);
not G2203 (W806, W2203);
not G2204 (W807, W2204);
not G2205 (W808, W2205);
not G2206 (W809, W2206);
not G2207 (W810, W2207);
not G2208 (W811, W2208);
not G2209 (W812, W2209);
not G2210 (W813, W2210);
not G2211 (W814, W2211);
not G2212 (W815, W2212);
not G2213 (W816, W2213);
not G2214 (W817, W2214);
not G2215 (W818, W2215);
not G2216 (W819, W2216);
not G2217 (W820, W2217);
not G2218 (W821, W2218);
not G2219 (W822, W2219);
not G2220 (W823, W2220);
not G2221 (W824, W2221);
not G2222 (W825, W2222);
not G2223 (W826, W2223);
not G2224 (W827, W2224);
not G2225 (W828, W2225);
not G2226 (W829, W2226);
not G2227 (W830, W2227);
not G2228 (W831, W2228);
not G2229 (W832, W2229);
not G2230 (W833, W2230);
not G2231 (W834, W2231);
not G2232 (W835, W2232);
not G2233 (W836, W2233);
not G2234 (W837, W2234);
not G2235 (W838, W2235);
not G2236 (W839, W2236);
not G2237 (W840, W2237);
not G2238 (W841, W2238);
not G2239 (W842, W2239);
not G2240 (W843, W2240);
not G2241 (W844, W2241);
not G2242 (W845, W2242);
not G2243 (W846, W2243);
not G2244 (W847, W2244);
not G2245 (W848, W2245);
not G2246 (W849, W2246);
not G2247 (W850, W2247);
not G2248 (W851, W2248);
not G2249 (W852, W2249);
not G2250 (W853, W2250);
not G2251 (W854, W2251);
not G2252 (W855, W2252);
not G2253 (W856, W2253);
not G2254 (W857, W2254);
not G2255 (W858, W2255);
not G2256 (W859, W2256);
not G2257 (W860, W2257);
not G2258 (W861, W2258);
not G2259 (W862, W2259);
not G2260 (W863, W2260);
not G2261 (W864, W2261);
not G2262 (W865, W2262);
not G2263 (W866, W2263);
not G2264 (W867, W2264);
not G2265 (W868, W2265);
not G2266 (W869, W2266);
not G2267 (W870, W2267);
not G2268 (W871, W2268);
not G2269 (W872, W2269);
not G2270 (W873, W2270);
not G2271 (W874, W2271);
not G2272 (W875, W2272);
not G2273 (W876, W2273);
not G2274 (W877, W2274);
not G2275 (W878, W2275);
not G2276 (W879, W2276);
not G2277 (W880, W2277);
not G2278 (W881, W2278);
not G2279 (W882, W2279);
not G2280 (W883, W2280);
not G2281 (W884, W2281);
not G2282 (W885, W2282);
not G2283 (W886, W2283);
not G2284 (W887, W2284);
not G2285 (W888, W2285);
not G2286 (W889, W2286);
not G2287 (W890, W2287);
not G2288 (W891, W2288);
not G2289 (W892, W2289);
not G2290 (W893, W2290);
not G2291 (W894, W2291);
not G2292 (W895, W2292);
not G2293 (W896, W2293);
not G2294 (W897, W2294);
not G2295 (W898, W2295);
not G2296 (W899, W2296);
not G2297 (W900, W2297);
not G2298 (W901, W2298);
not G2299 (W902, W2299);
not G2300 (W903, W2300);
not G2301 (W904, W2301);
not G2302 (W905, W2302);
not G2303 (W906, W2303);
not G2304 (W907, W2304);
not G2305 (W908, W2305);
not G2306 (W909, W2306);
not G2307 (W910, W2307);
not G2308 (W911, W2308);
not G2309 (W912, W2309);
not G2310 (W913, W2310);
not G2311 (W914, W2311);
not G2312 (W915, W2312);
not G2313 (W916, W2313);
not G2314 (W917, W2314);
not G2315 (W918, W2315);
not G2316 (W919, W2316);
not G2317 (W920, W2317);
not G2318 (W921, W2318);
not G2319 (W922, W2319);
not G2320 (W923, W2320);
not G2321 (W924, W2321);
not G2322 (W925, W2322);
not G2323 (W926, W2323);
not G2324 (W927, W2324);
not G2325 (W928, W2325);
not G2326 (W929, W2326);
not G2327 (W930, W2327);
not G2328 (W931, W2328);
not G2329 (W932, W2329);
not G2330 (W933, W2330);
not G2331 (W934, W2331);
not G2332 (W935, W2332);
not G2333 (W936, W2333);
not G2334 (W937, W2334);
not G2335 (W938, W2335);
not G2336 (W939, W2336);
not G2337 (W940, W2337);
not G2338 (W941, W2338);
not G2339 (W942, W2339);
not G2340 (W943, W2340);
not G2341 (W944, W2341);
not G2342 (W945, W2342);
not G2343 (W946, W2343);
not G2344 (W947, W2344);
not G2345 (W948, W2345);
not G2346 (W949, W2346);
not G2347 (W950, W2347);
not G2348 (W951, W2348);
not G2349 (W952, W2349);
not G2350 (W953, W2350);
not G2351 (W954, W2351);
not G2352 (W955, W2352);
not G2353 (W956, W2353);
not G2354 (W957, W2354);
not G2355 (W958, W2355);
not G2356 (W959, W2356);
not G2357 (W960, W2357);
not G2358 (W961, W2358);
not G2359 (W962, W2359);
not G2360 (W963, W2360);
not G2361 (W964, W2361);
not G2362 (W965, W2362);
not G2363 (W966, W2363);
not G2364 (W967, W2364);
not G2365 (W968, W2365);
not G2366 (W969, W2366);
not G2367 (W970, W2367);
not G2368 (W971, W2368);
not G2369 (W972, W2369);
not G2370 (W973, W2370);
not G2371 (W974, W2371);
not G2372 (W975, W2372);
not G2373 (W976, W2373);
not G2374 (W977, W2374);
not G2375 (W978, W2375);
not G2376 (W979, W2376);
not G2377 (W980, W2377);
not G2378 (W981, W2378);
not G2379 (W982, W2379);
not G2380 (W983, W2380);
not G2381 (W984, W2381);
not G2382 (W985, W2382);
not G2383 (W986, W2383);
not G2384 (W987, W2384);
not G2385 (W988, W2385);
not G2386 (W989, W2386);
not G2387 (W990, W2387);
not G2388 (W991, W2388);
not G2389 (W992, W2389);
not G2390 (W993, W2390);
not G2391 (W994, W2391);
not G2392 (W995, W2392);
not G2393 (W996, W2393);
not G2394 (W997, W2394);
not G2395 (W998, W2395);
not G2396 (W999, W2396);
not G2397 (W1000, W2397);
not G2398 (W1001, W2398);
not G2399 (W1002, W2399);
not G2400 (W1003, W2400);
not G2401 (W1004, W2401);
not G2402 (W1005, W2402);
not G2403 (W1006, W2403);
not G2404 (W1007, W2404);
not G2405 (W1008, W2405);
not G2406 (W1009, W2406);
not G2407 (W1010, W2407);
not G2408 (W1011, W2408);
not G2409 (W1012, W2409);
not G2410 (W1013, W2410);
not G2411 (W1014, W2411);
not G2412 (W1015, W2412);
not G2413 (W1016, W2413);
not G2414 (W1017, W2414);
not G2415 (W1018, W2415);
not G2416 (W1019, W2416);
not G2417 (W1020, W2417);
not G2418 (W1021, W2418);
not G2419 (W1022, W2419);
not G2420 (W1023, W2420);
not G2421 (W1024, W2421);
not G2422 (W1025, W2422);
not G2423 (W1026, W2423);
not G2424 (W1027, W2424);
not G2425 (W1028, W2425);
not G2426 (W1029, W2426);
not G2427 (W1030, W2427);
not G2428 (W1031, W2428);
not G2429 (W1032, W2429);
not G2430 (W1033, W2430);
not G2431 (W1034, W2431);
not G2432 (W1035, W2432);
not G2433 (W1036, W2433);
not G2434 (W1037, W2434);
not G2435 (W1038, W2435);
not G2436 (W1039, W2436);
not G2437 (W1040, W2437);
not G2438 (W1041, W2438);
not G2439 (W1042, W2439);
not G2440 (W1043, W2440);
not G2441 (W1044, W2441);
not G2442 (W1045, W2442);
not G2443 (W1046, W2443);
not G2444 (W1047, W2444);
not G2445 (W1048, W2445);
not G2446 (W1049, W2446);
not G2447 (W1050, W2447);
not G2448 (W1051, W2448);
not G2449 (W1052, W2449);
not G2450 (W1053, W2450);
not G2451 (W1054, W2451);
not G2452 (W1055, W2452);
not G2453 (W1056, W2453);
not G2454 (W1057, W2454);
not G2455 (W1058, W2455);
not G2456 (W1059, W2456);
not G2457 (W1060, W2457);
not G2458 (W1061, W2458);
not G2459 (W1062, W2459);
not G2460 (W1063, W2460);
not G2461 (W1064, W2461);
not G2462 (W1065, W2462);
not G2463 (W1066, W2463);
not G2464 (W1067, W2464);
not G2465 (W1068, W2465);
not G2466 (W1069, W2466);
not G2467 (W1070, W2467);
not G2468 (W1071, W2468);
not G2469 (W1072, W2469);
not G2470 (W1073, W2470);
not G2471 (W1074, W2471);
not G2472 (W1075, W2472);
not G2473 (W1076, W2473);
not G2474 (W1077, W2474);
not G2475 (W1078, W2475);
not G2476 (W1079, W2476);
not G2477 (W1080, W2477);
not G2478 (W1081, W2478);
not G2479 (W1082, W2479);
not G2480 (W1083, W2480);
not G2481 (W1084, W2481);
not G2482 (W1085, W2482);
not G2483 (W1086, W2483);
not G2484 (W1087, W2484);
not G2485 (W1088, W2485);
not G2486 (W1089, W2486);
not G2487 (W1090, W2487);
not G2488 (W1091, W2488);
not G2489 (W1092, W2489);
not G2490 (W1093, W2490);
not G2491 (W1094, W2491);
not G2492 (W1095, W2492);
not G2493 (W1096, W2493);
not G2494 (W1097, W2494);
not G2495 (W1098, W2495);
not G2496 (W1099, W2496);
not G2497 (W1100, W2497);
not G2498 (W1101, W2498);
not G2499 (W1102, W2499);
not G2500 (W1103, W2500);
not G2501 (W1104, W2501);
not G2502 (W1105, W2502);
not G2503 (W1106, W2503);
not G2504 (W1107, W2504);
not G2505 (W1108, W2505);
not G2506 (W1109, W2506);
not G2507 (W1110, W2507);
not G2508 (W1111, W2508);
not G2509 (W1112, W2509);
not G2510 (W1113, W2510);
not G2511 (W1114, W2511);
not G2512 (W1115, W2512);
not G2513 (W1116, W2513);
not G2514 (W1117, W2514);
not G2515 (W1118, W2515);
not G2516 (W1119, W2516);
not G2517 (W1120, W2517);
not G2518 (W1121, W2518);
not G2519 (W1122, W2519);
not G2520 (W1123, W2520);
not G2521 (W1124, W2521);
not G2522 (W1125, W2522);
not G2523 (W1126, W2523);
not G2524 (W1127, W2524);
not G2525 (W1128, W2525);
not G2526 (W1129, W2526);
not G2527 (W1130, W2527);
not G2528 (W1131, W2528);
not G2529 (W1132, W2529);
not G2530 (W1133, W2530);
not G2531 (W1134, W2531);
not G2532 (W1135, W2532);
not G2533 (W1136, W2533);
not G2534 (W1137, W2534);
not G2535 (W1138, W2535);
not G2536 (W1139, W2536);
not G2537 (W1140, W2537);
not G2538 (W1141, W2538);
not G2539 (W1142, W2539);
not G2540 (W1143, W2540);
not G2541 (W1144, W2541);
not G2542 (W1145, W2542);
not G2543 (W1146, W2543);
not G2544 (W1147, W2544);
not G2545 (W1148, W2545);
not G2546 (W1149, W2546);
not G2547 (W1150, W2547);
not G2548 (W1151, W2548);
not G2549 (W1152, W2549);
not G2550 (W1153, W2550);
not G2551 (W1154, W2551);
not G2552 (W1155, W2552);
not G2553 (W1156, W2553);
not G2554 (W1157, W2554);
not G2555 (W1158, W2555);
not G2556 (W1159, W2556);
not G2557 (W1160, W2557);
not G2558 (W1161, W2558);
not G2559 (W1162, W2559);
not G2560 (W1163, W2560);
not G2561 (W1164, W2561);
not G2562 (W1165, W2562);
not G2563 (W1166, W2563);
not G2564 (W1167, W2564);
not G2565 (W1168, W2565);
not G2566 (W1169, W2566);
not G2567 (W1170, W2567);
not G2568 (W1171, W2568);
not G2569 (W1172, W2569);
not G2570 (W1173, W2570);
not G2571 (W1174, W2571);
not G2572 (W1175, W2572);
not G2573 (W1176, W2573);
not G2574 (W1177, W2574);
not G2575 (W1178, W2575);
not G2576 (W1179, W2576);
not G2577 (W1180, W2577);
not G2578 (W1181, W2578);
not G2579 (W1182, W2579);
not G2580 (W1183, W2580);
not G2581 (W1184, W2581);
not G2582 (W1185, W2582);
not G2583 (W1186, W2583);
not G2584 (W1187, W2584);
not G2585 (W1188, W2585);
not G2586 (W1189, W2586);
not G2587 (W1190, W2587);
not G2588 (W1191, W2588);
not G2589 (W1192, W2589);
not G2590 (W1193, W2590);
not G2591 (W1194, W2591);
not G2592 (W1195, W2592);
not G2593 (W1196, W2593);
not G2594 (W1197, W2594);
not G2595 (W1198, W2595);
not G2596 (W1199, W2596);
not G2597 (W1200, W2597);
not G2598 (W1201, W2598);
not G2599 (W1202, W2599);
not G2600 (W1203, W2600);
not G2601 (W1204, W2601);
not G2602 (W1205, W2602);
not G2603 (W1206, W2603);
not G2604 (W1207, W2604);
not G2605 (W1208, W2605);
not G2606 (W1209, W2606);
not G2607 (W1210, W2607);
not G2608 (W1211, W2608);
not G2609 (W1212, W2609);
not G2610 (W1213, W2610);
not G2611 (W1214, W2611);
not G2612 (W1215, W2612);
not G2613 (W1216, W2613);
not G2614 (W1217, W2614);
not G2615 (W1218, W2615);
not G2616 (W1219, W2616);
not G2617 (W1220, W2617);
not G2618 (W1221, W2618);
not G2619 (W1222, W2619);
not G2620 (W1223, W2620);
not G2621 (W1224, W2621);
not G2622 (W1225, W2622);
not G2623 (W1226, W2623);
not G2624 (W1227, W2624);
not G2625 (W1228, W2625);
not G2626 (W1229, W2626);
not G2627 (W1230, W2627);
not G2628 (W1231, W2628);
not G2629 (W1232, W2629);
not G2630 (W1233, W2630);
not G2631 (W1234, W2631);
not G2632 (W1235, W2632);
not G2633 (W1236, W2633);
not G2634 (W1237, W2634);
not G2635 (W1238, W2635);
not G2636 (W1239, W2636);
not G2637 (W1240, W2637);
not G2638 (W1241, W2638);
not G2639 (W1242, W2639);
not G2640 (W1243, W2640);
not G2641 (W1244, W2641);
not G2642 (W1245, W2642);
not G2643 (W1246, W2643);
not G2644 (W1247, W2644);
not G2645 (W1248, W2645);
not G2646 (W1249, W2646);
not G2647 (W1250, W2647);
not G2648 (W1251, W2648);
not G2649 (W1252, W2649);
not G2650 (W1253, W2650);
not G2651 (W1254, W2651);
not G2652 (W1255, W2652);
not G2653 (W1256, W2653);
not G2654 (W1257, W2654);
not G2655 (W1258, W2655);
not G2656 (W1259, W2656);
not G2657 (W1260, W2657);
not G2658 (W1261, W2658);
not G2659 (W1262, W2659);
not G2660 (W1263, W2660);
not G2661 (W1264, W2661);
not G2662 (W1265, W2662);
not G2663 (W1266, W2663);
not G2664 (W1267, W2664);
not G2665 (W1268, W2665);
not G2666 (W1269, W2666);
not G2667 (W1270, W2667);
not G2668 (W1271, W2668);
not G2669 (W1272, W2669);
not G2670 (W1273, W2670);
not G2671 (W1274, W2671);
not G2672 (W1275, W2672);
not G2673 (W1276, W2673);
not G2674 (W1277, W2674);
not G2675 (W1278, W2675);
not G2676 (W1279, W2676);
not G2677 (W1280, W2677);
not G2678 (W1281, W2678);
not G2679 (W1282, W2679);
not G2680 (W1283, W2680);
not G2681 (W1284, W2681);
not G2682 (W1285, W2682);
not G2683 (W1286, W2683);
not G2684 (W1287, W2684);
not G2685 (W1288, W2685);
not G2686 (W1289, W2686);
not G2687 (W1290, W2687);
not G2688 (W1291, W2688);
not G2689 (W1292, W2689);
not G2690 (W1293, W2690);
not G2691 (W1294, W2691);
not G2692 (W1295, W2692);
not G2693 (W1296, W2693);
not G2694 (W1297, W2694);
not G2695 (W1298, W2695);
not G2696 (W1299, W2696);
not G2697 (W1300, W2697);
not G2698 (W1301, W2698);
not G2699 (W1302, W2699);
not G2700 (W1303, W2700);
not G2701 (W1304, W2701);
not G2702 (W1305, W2702);
not G2703 (W1306, W2703);
not G2704 (W1307, W2704);
not G2705 (W1308, W2705);
not G2706 (W1309, W2706);
not G2707 (W1310, W2707);
not G2708 (W1311, W2708);
not G2709 (W1312, W2709);
not G2710 (W1313, W2710);
not G2711 (W1314, W2711);
not G2712 (W1315, W2712);
not G2713 (W1316, W2713);
not G2714 (W1317, W2714);
not G2715 (W1318, W2715);
not G2716 (W1319, W2716);
not G2717 (W1320, W2717);
not G2718 (W1321, W2718);
not G2719 (W1322, W2719);
not G2720 (W1323, W2720);
not G2721 (W1324, W2721);
not G2722 (W1325, W2722);
not G2723 (W1326, W2723);
not G2724 (W1327, W2724);
not G2725 (W1328, W2725);
not G2726 (W1329, W2726);
not G2727 (W1330, W2727);
not G2728 (W1331, W2728);
not G2729 (W1332, W2729);
not G2730 (W1333, W2730);
not G2731 (W1334, W2731);
not G2732 (W1335, W2732);
not G2733 (W1336, W2733);
not G2734 (W1337, W2734);
not G2735 (W1338, W2735);
not G2736 (W1339, W2736);
not G2737 (W1340, W2737);
not G2738 (W1341, W2738);
not G2739 (W1342, W2739);
not G2740 (W1343, W2740);
not G2741 (W1344, W2741);
not G2742 (W1345, W2742);
not G2743 (W1346, W2743);
not G2744 (W1347, W2744);
not G2745 (W1348, W2745);
not G2746 (W1349, W2746);
not G2747 (W1350, W2747);
not G2748 (W1351, W2748);
not G2749 (W1352, W2749);
not G2750 (W1353, W2750);
not G2751 (W1354, W2751);
not G2752 (W1355, W2752);
not G2753 (W1356, W2753);
not G2754 (W1357, W2754);
not G2755 (W1358, W2755);
not G2756 (W1359, W2756);
not G2757 (W1360, W2757);
not G2758 (W1361, W2758);
not G2759 (W1362, W2759);
not G2760 (W1363, W2760);
not G2761 (W1364, W2761);
not G2762 (W1365, W2762);
not G2763 (W1366, W2763);
not G2764 (W1367, W2764);
not G2765 (W1368, W2765);
not G2766 (W1369, W2766);
not G2767 (W1370, W2767);
not G2768 (W1371, W2768);
not G2769 (W1372, W2769);
not G2770 (W1373, W2770);
not G2771 (W1374, W2771);
not G2772 (W1375, W2772);
not G2773 (W1376, W2773);
not G2774 (W1377, W2774);
not G2775 (W1378, W2775);
not G2776 (W1379, W2776);
not G2777 (W1380, W2777);
not G2778 (W1381, W2778);
not G2779 (W1382, W2779);
not G2780 (W1383, W2780);
not G2781 (W1384, W2781);
not G2782 (W1385, W2782);
not G2783 (W1386, W2783);
not G2784 (W1387, W2784);
not G2785 (W1388, W2785);
not G2786 (W1389, W2786);
not G2787 (W1390, W2787);
not G2788 (W1391, W2788);
not G2789 (W1392, W2789);
not G2790 (W1393, W2790);
not G2791 (W1394, W2791);
not G2792 (W1395, W2792);
not G2793 (W1396, W2793);
not G2794 (W1397, W2794);
not G2795 (W1398, W2795);
not G2796 (W1399, W2796);
not G2797 (W1400, W2797);
not G2798 (W1401, W2798);
not G2799 (W1402, W2799);
not G2800 (W1403, W2800);
not G2801 (W1404, W2801);
not G2802 (W1405, W2802);
not G2803 (W1406, W2803);
not G2804 (W1407, W2804);
not G2805 (W1408, W2805);
not G2806 (W1409, W2806);
not G2807 (W1410, W2807);
not G2808 (W1411, W2808);
not G2809 (W1412, W2809);
not G2810 (W1413, W2810);
not G2811 (W1414, W2811);
not G2812 (W1415, W2812);
not G2813 (W1416, W2813);
not G2814 (W1417, W2814);
not G2815 (W1418, W2815);
not G2816 (W1419, W2816);
not G2817 (W1420, W2817);
not G2818 (W1421, W2818);
not G2819 (W1422, W2819);
not G2820 (W1423, W2820);
not G2821 (W1424, W2821);
not G2822 (W1425, W2822);
not G2823 (W1426, W2823);
not G2824 (W1427, W2824);
not G2825 (W1428, W2825);
not G2826 (W1429, W2826);
not G2827 (W1430, W2827);
not G2828 (W1431, W2828);
not G2829 (W1432, W2829);
not G2830 (W1433, W2830);
not G2831 (W1434, W2831);
not G2832 (W1435, W2832);
not G2833 (W1436, W2833);
not G2834 (W1437, W2834);
not G2835 (W1438, W2835);
not G2836 (W1439, W2836);
not G2837 (W1440, W2837);
not G2838 (W1441, W2838);
not G2839 (W1442, W2839);
not G2840 (W1443, W2840);
not G2841 (W1444, W2841);
not G2842 (W1445, W2842);
not G2843 (W1446, W2843);
not G2844 (W1447, W2844);
not G2845 (W1448, W2845);
not G2846 (W1449, W2846);
not G2847 (W1450, W2847);
not G2848 (W1451, W2848);
not G2849 (W1452, W2849);
not G2850 (W1453, W2850);
not G2851 (W1454, W2851);
not G2852 (W1455, W2852);
not G2853 (W1456, W2853);
not G2854 (W1457, W2854);
not G2855 (W1458, W2855);
not G2856 (W1459, W2856);
not G2857 (W1460, W2857);
not G2858 (W1461, W2858);
not G2859 (W1462, W2859);
not G2860 (W1463, W2860);
not G2861 (W1464, W2861);
not G2862 (W1465, W2862);
not G2863 (W1466, W2863);
not G2864 (W1467, W2864);
not G2865 (W1468, W2865);
not G2866 (W1469, W2866);
not G2867 (W1470, W2867);
not G2868 (W1471, W2868);
not G2869 (W1472, W2869);
not G2870 (W1473, W2870);
not G2871 (W1474, W2871);
not G2872 (W1475, W2872);
not G2873 (W1476, W2873);
not G2874 (W1477, W2874);
not G2875 (W1478, W2875);
not G2876 (W1479, W2876);
not G2877 (W1480, W2877);
not G2878 (W1481, W2878);
not G2879 (W1482, W2879);
not G2880 (W1483, W2880);
not G2881 (W1484, W2881);
not G2882 (W1485, W2882);
not G2883 (W1486, W2883);
not G2884 (W1487, W2884);
not G2885 (W1488, W2885);
not G2886 (W1489, W2886);
not G2887 (W1490, W2887);
not G2888 (W1491, W2888);
not G2889 (W1492, W2889);
not G2890 (W1493, W2890);
not G2891 (W1494, W2891);
not G2892 (W1495, W2892);
not G2893 (W1496, W2893);
not G2894 (W1497, W2894);
not G2895 (W1498, W2895);
not G2896 (W1499, W2896);
not G2897 (W1500, W2897);
not G2898 (W1501, W2898);
not G2899 (W1502, W2899);
not G2900 (W1503, W2900);
not G2901 (W1504, W2901);
not G2902 (W1505, W2902);
not G2903 (W1506, W2903);
not G2904 (W1507, W2904);
not G2905 (W1508, W2905);
not G2906 (W1509, W2906);
not G2907 (W1510, W2907);
not G2908 (W1511, W2908);
not G2909 (W1512, W2909);
not G2910 (W1513, W2910);
not G2911 (W1514, W2911);
not G2912 (W1515, W2912);
not G2913 (W1516, W2913);
not G2914 (W1517, W2914);
not G2915 (W1518, W2915);
not G2916 (W1519, W2916);
not G2917 (W1520, W2917);
not G2918 (W1521, W2918);
not G2919 (W1522, W2919);
not G2920 (W1523, W2920);
not G2921 (W1524, W2921);
not G2922 (W1525, W2922);
not G2923 (W1526, W2923);
not G2924 (W1527, W2924);
not G2925 (W1528, W2925);
not G2926 (W1529, W2926);
not G2927 (W1530, W2927);
not G2928 (W1531, W2928);
not G2929 (W1532, W2929);
not G2930 (W1533, W2930);
not G2931 (W1534, W2931);
not G2932 (W1535, W2932);
not G2933 (W1536, W2933);
not G2934 (W1537, W2934);
not G2935 (W1538, W2935);
not G2936 (W1539, W2936);
not G2937 (W1540, W2937);
not G2938 (W1541, W2938);
not G2939 (W1542, W2939);
not G2940 (W1543, W2940);
not G2941 (W1544, W2941);
not G2942 (W1545, W2942);
not G2943 (W1546, W2943);
not G2944 (W1547, W2944);
not G2945 (W1548, W2945);
not G2946 (W1549, W2946);
not G2947 (W1550, W2947);
not G2948 (W1551, W2948);
not G2949 (W1552, W2949);
not G2950 (W1553, W2950);
not G2951 (W1554, W2951);
not G2952 (W1555, W2952);
not G2953 (W1556, W2953);
not G2954 (W1557, W2954);
not G2955 (W1558, W2955);
not G2956 (W1559, W2956);
not G2957 (W1560, W2957);
not G2958 (W1561, W2958);
not G2959 (W1562, W2959);
not G2960 (W1563, W2960);
not G2961 (W1564, W2961);
not G2962 (W1565, W2962);
not G2963 (W1566, W2963);
not G2964 (W1567, W2964);
not G2965 (W1568, W2965);
not G2966 (W1569, W2966);
not G2967 (W1570, W2967);
not G2968 (W1571, W2968);
not G2969 (W1572, W2969);
not G2970 (W1573, W2970);
not G2971 (W1574, W2971);
not G2972 (W1575, W2972);
not G2973 (W1576, W2973);
not G2974 (W1577, W2974);
not G2975 (W1578, W2975);
not G2976 (W1579, W2976);
not G2977 (W1580, W2977);
not G2978 (W1581, W2978);
not G2979 (W1582, W2979);
not G2980 (W1583, W2980);
not G2981 (W1584, W2981);
not G2982 (W1585, W2982);
not G2983 (W1586, W2983);
not G2984 (W1587, W2984);
not G2985 (W1588, W2985);
not G2986 (W1589, W2986);
not G2987 (W1590, W2987);
not G2988 (W1591, W2988);
not G2989 (W1592, W2989);
not G2990 (W1593, W2990);
not G2991 (W1594, W2991);
not G2992 (W1595, W2992);
not G2993 (W1596, W2993);
not G2994 (W1597, W2994);
not G2995 (W1598, W2995);
not G2996 (W1599, W2996);
not G2997 (W1600, W2997);
not G2998 (W1601, W2998);
not G2999 (W1602, W2999);
not G3000 (W1603, W3000);
not G3001 (W1604, W3001);
not G3002 (W1605, W3002);
not G3003 (W1606, W3003);
not G3004 (W1607, W3004);
not G3005 (W1608, W3005);
not G3006 (W1609, W3006);
not G3007 (W1610, W3007);
not G3008 (W1611, W3008);
not G3009 (W1612, W3009);
not G3010 (W1613, W3010);
not G3011 (W1614, W3011);
not G3012 (W1615, W3012);
not G3013 (W1616, W3013);
not G3014 (W1617, W3014);
not G3015 (W1618, W3015);
not G3016 (W1619, W3016);
not G3017 (W1620, W3017);
not G3018 (W1621, W3018);
not G3019 (W1622, W3019);
not G3020 (W1623, W3020);
not G3021 (W1624, W3021);
not G3022 (W1625, W3022);
not G3023 (W1626, W3023);
not G3024 (W1627, W3024);
not G3025 (W1628, W3025);
not G3026 (W1629, W3026);
not G3027 (W1630, W3027);
not G3028 (W1631, W3028);
not G3029 (W1632, W3029);
not G3030 (W1633, W3030);
not G3031 (W1634, W3031);
not G3032 (W1635, W3032);
not G3033 (W1636, W3033);
not G3034 (W1637, W3034);
not G3035 (W1638, W3035);
not G3036 (W1639, W3036);
not G3037 (W1640, W3037);
not G3038 (W1641, W3038);
not G3039 (W1642, W3039);
not G3040 (W1643, W3040);
not G3041 (W1644, W3041);
not G3042 (W1645, W3042);
not G3043 (W1646, W3043);
not G3044 (W1647, W3044);
not G3045 (W1648, W3045);
not G3046 (W1649, W3046);
not G3047 (W1650, W3047);
not G3048 (W1651, W3048);
not G3049 (W1652, W3049);
not G3050 (W1653, W3050);
not G3051 (W1654, W3051);
not G3052 (W1655, W3052);
not G3053 (W1656, W3053);
not G3054 (W1657, W3054);
not G3055 (W1658, W3055);
not G3056 (W1659, W3056);
not G3057 (W1660, W3057);
not G3058 (W1661, W3058);
not G3059 (W1662, W3059);
not G3060 (W1663, W3060);
not G3061 (W1664, W3061);
not G3062 (W1665, W3062);
not G3063 (W1666, W3063);
not G3064 (W1667, W3064);
not G3065 (W1668, W3065);
not G3066 (W1669, W3066);
not G3067 (W1670, W3067);
not G3068 (W1671, W3068);
not G3069 (W1672, W3069);
not G3070 (W1673, W3070);
not G3071 (W1674, W3071);
not G3072 (W1675, W3072);
not G3073 (W1676, W3073);
not G3074 (W1677, W3074);
not G3075 (W1678, W3075);
not G3076 (W1679, W3076);
not G3077 (W1680, W3077);
not G3078 (W1681, W3078);
not G3079 (W1682, W3079);
not G3080 (W1683, W3080);
not G3081 (W1684, W3081);
not G3082 (W1685, W3082);
not G3083 (W1686, W3083);
not G3084 (W1687, W3084);
not G3085 (W1688, W3085);
not G3086 (W1689, W3086);
not G3087 (W1690, W3087);
not G3088 (W1691, W3088);
not G3089 (W1692, W3089);
not G3090 (W1693, W3090);
not G3091 (W1694, W3091);
not G3092 (W1695, W3092);
not G3093 (W1696, W3093);
not G3094 (W1697, W3094);
not G3095 (W1698, W3095);
not G3096 (W1699, W3096);
not G3097 (W1700, W3097);
not G3098 (W1701, W3098);
not G3099 (W1702, W3099);
not G3100 (W1703, W3100);
not G3101 (W1704, W3101);
not G3102 (W1705, W3102);
not G3103 (W1706, W3103);
not G3104 (W1707, W3104);
not G3105 (W1708, W3105);
not G3106 (W1709, W3106);
not G3107 (W1710, W3107);
not G3108 (W1711, W3108);
not G3109 (W1712, W3109);
not G3110 (W1713, W3110);
not G3111 (W1714, W3111);
not G3112 (W1715, W3112);
not G3113 (W1716, W3113);
not G3114 (W1717, W3114);
not G3115 (W1718, W3115);
not G3116 (W1719, W3116);
not G3117 (W1720, W3117);
not G3118 (W1721, W3118);
not G3119 (W1722, W3119);
not G3120 (W1723, W3120);
not G3121 (W1724, W3121);
not G3122 (W1725, W3122);
not G3123 (W1726, W3123);
not G3124 (W1727, W3124);
not G3125 (W1728, W3125);
not G3126 (W1729, W3126);
not G3127 (W1730, W3127);
not G3128 (W1731, W3128);
not G3129 (W1732, W3129);
not G3130 (W1733, W3130);
not G3131 (W1734, W3131);
not G3132 (W1735, W3132);
not G3133 (W1736, W3133);
not G3134 (W1737, W3134);
not G3135 (W1738, W3135);
not G3136 (W1739, W3136);
not G3137 (W1740, W3137);
not G3138 (W1741, W3138);
not G3139 (W1742, W3139);
not G3140 (W1743, W3140);
not G3141 (W1744, W3141);
not G3142 (W1745, W3142);
not G3143 (W1746, W3143);
not G3144 (W1747, W3144);
not G3145 (W1748, W3145);
not G3146 (W1749, W3146);
not G3147 (W1750, W3147);
not G3148 (W1751, W3148);
not G3149 (W1752, W3149);
not G3150 (W1753, W3150);
not G3151 (W1754, W3151);
not G3152 (W1755, W3152);
not G3153 (W1756, W3153);
not G3154 (W1757, W3154);
not G3155 (W1758, W3155);
not G3156 (W1759, W3156);
not G3157 (W1760, W3157);
not G3158 (W1761, W3158);
not G3159 (W1762, W3159);
not G3160 (W1763, W3160);
not G3161 (W1764, W3161);
not G3162 (W1765, W3162);
not G3163 (W1766, W3163);
not G3164 (W1767, W3164);
not G3165 (W1768, W3165);
not G3166 (W1769, W3166);
not G3167 (W1770, W3167);
not G3168 (W1771, W3168);
not G3169 (W1772, W3169);
not G3170 (W1773, W3170);
not G3171 (W1774, W3171);
not G3172 (W1775, W3172);
not G3173 (W1776, W3173);
not G3174 (W1777, W3174);
not G3175 (W1778, W3175);
not G3176 (W1779, W3176);
not G3177 (W1780, W3177);
not G3178 (W1781, W3178);
not G3179 (W1782, W3179);
not G3180 (W1783, W3180);
not G3181 (W1784, W3181);
not G3182 (W1785, W3182);
not G3183 (W1786, W3183);
not G3184 (W1787, W3184);
not G3185 (W1788, W3185);
not G3186 (W1789, W3186);
not G3187 (W1790, W3187);
not G3188 (W1791, W3188);
not G3189 (W1792, W3189);
not G3190 (W1793, W3190);
not G3191 (W1794, W3191);
not G3192 (W1795, W3192);
not G3193 (W1796, W3193);
not G3194 (W1797, W3194);
not G3195 (W1798, W3195);
not G3196 (W1799, W3196);
not G3197 (W1800, W3197);
not G3198 (W1801, W3198);
not G3199 (W1802, W3199);
not G3200 (W1803, W3200);
not G3201 (W1804, W3201);
not G3202 (W1805, W3202);
not G3203 (W1806, W3203);
not G3204 (W1807, W3204);
not G3205 (W1808, W3205);
not G3206 (W1809, W3206);
not G3207 (W1810, W3207);
not G3208 (W1811, W3208);
not G3209 (W1812, W3209);
not G3210 (W1813, W3210);
not G3211 (W1814, W3211);
not G3212 (W1815, W3212);
not G3213 (W1816, W3213);
not G3214 (W1817, W3214);
not G3215 (W1818, W3215);
not G3216 (W1819, W3216);
not G3217 (W1820, W3217);
not G3218 (W1821, W3218);
not G3219 (W1822, W3219);
not G3220 (W1823, W3220);
not G3221 (W1824, W3221);
not G3222 (W1825, W3222);
not G3223 (W1826, W3223);
not G3224 (W1827, W3224);
not G3225 (W1828, W3225);
not G3226 (W1829, W3226);
not G3227 (W1830, W3227);
not G3228 (W1831, W3228);
not G3229 (W1832, W3229);
not G3230 (W1833, W3230);
not G3231 (W1834, W3231);
not G3232 (W1835, W3232);
not G3233 (W1836, W3233);
not G3234 (W1837, W3234);
not G3235 (W1838, W3235);
not G3236 (W1839, W3236);
not G3237 (W1840, W3237);
not G3238 (W1841, W3238);
not G3239 (W1842, W3239);
not G3240 (W1843, W3240);
not G3241 (W1844, W3241);
not G3242 (W1845, W3242);
not G3243 (W1846, W3243);
not G3244 (W1847, W3244);
not G3245 (W1848, W3245);
not G3246 (W1849, W3246);
not G3247 (W1850, W3247);
not G3248 (W1851, W3248);
not G3249 (W1852, W3249);
not G3250 (W1853, W3250);
not G3251 (W1854, W3251);
not G3252 (W1855, W3252);
not G3253 (W1856, W3253);
not G3254 (W1857, W3254);
not G3255 (W1858, W3255);
not G3256 (W1859, W3256);
not G3257 (W1860, W3257);
not G3258 (W1861, W3258);
not G3259 (W1862, W3259);
not G3260 (W1863, W3260);
not G3261 (W1864, W3261);
not G3262 (W1865, W3262);
not G3263 (W1866, W3263);
not G3264 (W1867, W3264);
not G3265 (W1868, W3265);
not G3266 (W1869, W3266);
not G3267 (W1870, W3267);
not G3268 (W1871, W3268);
not G3269 (W1872, W3269);
not G3270 (W1873, W3270);
not G3271 (W1874, W3271);
not G3272 (W1875, W3272);
not G3273 (W1876, W3273);
not G3274 (W1877, W3274);
not G3275 (W1878, W3275);
not G3276 (W1879, W3276);
not G3277 (W1880, W3277);
not G3278 (W1881, W3278);
not G3279 (W1882, W3279);
not G3280 (W1883, W3280);
not G3281 (W1884, W3281);
not G3282 (W1885, W3282);
not G3283 (W1886, W3283);
not G3284 (W1887, W3284);
not G3285 (W1888, W3285);
not G3286 (W1889, W3286);
not G3287 (W1890, W3287);
not G3288 (W1891, W3288);
not G3289 (W1892, W3289);
not G3290 (W1893, W3290);
not G3291 (W1894, W3291);
not G3292 (W1895, W3292);
not G3293 (W1896, W3293);
not G3294 (W1897, W3294);
not G3295 (W1898, W3295);
not G3296 (W1899, W3296);
not G3297 (W1900, W3297);
not G3298 (W1901, W3298);
not G3299 (W1902, W3299);
not G3300 (W1903, W3300);
not G3301 (W1904, W3301);
not G3302 (W1905, W3302);
not G3303 (W1906, W3303);
not G3304 (W1907, W3304);
not G3305 (W1908, W3305);
not G3306 (W1909, W3306);
not G3307 (W1910, W3307);
not G3308 (W1911, W3308);
not G3309 (W1912, W3309);
not G3310 (W1913, W3310);
not G3311 (W1914, W3311);
not G3312 (W1915, W3312);
not G3313 (W1916, W3313);
not G3314 (W1917, W3314);
not G3315 (W1918, W3315);
not G3316 (W1919, W3316);
not G3317 (W1920, W3317);
not G3318 (W1921, W3318);
not G3319 (W1922, W3319);
not G3320 (W1923, W3320);
not G3321 (W1924, W3321);
not G3322 (W1925, W3322);
not G3323 (W1926, W3323);
not G3324 (W1927, W3324);
not G3325 (W1928, W3325);
not G3326 (W1929, W3326);
not G3327 (W1930, W3327);
not G3328 (W1931, W3328);
not G3329 (W1932, W3329);
not G3330 (W1933, W3330);
not G3331 (W1934, W3331);
not G3332 (W1935, W3332);
not G3333 (W1936, W3333);
not G3334 (W1937, W3334);
not G3335 (W1938, W3335);
not G3336 (W1939, W3336);
not G3337 (W1940, W3337);
not G3338 (W1941, W3338);
not G3339 (W1942, W3339);
not G3340 (W1943, W3340);
not G3341 (W1944, W3341);
not G3342 (W1945, W3342);
not G3343 (W1946, W3343);
not G3344 (W1947, W3344);
not G3345 (W1948, W3345);
not G3346 (W1949, W3346);
not G3347 (W1950, W3347);
not G3348 (W1951, W3348);
not G3349 (W1952, W3349);
not G3350 (W1953, W3350);
not G3351 (W1954, W3351);
not G3352 (W1955, W3352);
not G3353 (W1956, W3353);
not G3354 (W1957, W3354);
not G3355 (W1958, W3355);
not G3356 (W1959, W3356);
not G3357 (W1960, W3357);
not G3358 (W1961, W3358);
not G3359 (W1962, W3359);
not G3360 (W1963, W3360);
not G3361 (W1964, W3361);
not G3362 (W1965, W3362);
not G3363 (W1966, W3363);
not G3364 (W1967, W3364);
not G3365 (W1968, W3365);
not G3366 (W1969, W3366);
not G3367 (W1970, W3367);
not G3368 (W1971, W3368);
not G3369 (W1972, W3369);
not G3370 (W1973, W3370);
not G3371 (W1974, W3371);
not G3372 (W1975, W3372);
not G3373 (W1976, W3373);
not G3374 (W1977, W3374);
not G3375 (W1978, W3375);
not G3376 (W1979, W3376);
not G3377 (W1980, W3377);
not G3378 (W1981, W3378);
not G3379 (W1982, W3379);
not G3380 (W1983, W3380);
not G3381 (W1984, W3381);
not G3382 (W1985, W3382);
not G3383 (W1986, W3383);
not G3384 (W1987, W3384);
not G3385 (W1988, W3385);
not G3386 (W1989, W3386);
not G3387 (W1990, W3387);
not G3388 (W1991, W3388);
not G3389 (W1992, W3389);
not G3390 (W1993, W3390);
not G3391 (W1994, W3391);
not G3392 (W1995, W3392);
not G3393 (W1996, W3393);
not G3394 (W1997, W3394);
not G3395 (W1998, W3395);
not G3396 (W1999, W3396);
not G3397 (W2000, W3397);
not G3398 (W2001, W3398);
not G3399 (W2002, W3399);
not G3400 (W2003, W3400);
not G3401 (W2004, W3401);
not G3402 (W2005, W3402);
not G3403 (W2006, W3403);
not G3404 (W2007, W3404);
not G3405 (W2008, W3405);
not G3406 (W2009, W3406);
not G3407 (W2010, W3407);
not G3408 (W2011, W3408);
not G3409 (W2012, W3409);
not G3410 (W2013, W3410);
not G3411 (W2014, W3411);
not G3412 (W2015, W3412);
not G3413 (W2016, W3413);
not G3414 (W2017, W3414);
not G3415 (W2018, W3415);
not G3416 (W2019, W3416);
not G3417 (W2020, W3417);
not G3418 (W2021, W3418);
not G3419 (W2022, W3419);
not G3420 (W2023, W3420);
not G3421 (W2024, W3421);
not G3422 (W2025, W3422);
not G3423 (W2026, W3423);
not G3424 (W2027, W3424);
not G3425 (W2028, W3425);
not G3426 (W2029, W3426);
not G3427 (W2030, W3427);
not G3428 (W2031, W3428);
not G3429 (W2032, W3429);
not G3430 (W2033, W3430);
not G3431 (W2034, W3431);
not G3432 (W2035, W3432);
not G3433 (W2036, W3433);
not G3434 (W2037, W3434);
not G3435 (W2038, W3435);
not G3436 (W2039, W3436);
not G3437 (W2040, W3437);
not G3438 (W2041, W3438);
not G3439 (W2042, W3439);
not G3440 (W2043, W3440);
not G3441 (W2044, W3441);
not G3442 (W2045, W3442);
not G3443 (W2046, W3443);
not G3444 (W2047, W3444);
not G3445 (W2048, W3445);
not G3446 (W2049, W3446);
not G3447 (W2050, W3447);
not G3448 (W2051, W3448);
not G3449 (W2052, W3449);
not G3450 (W2053, W3450);
not G3451 (W2054, W3451);
not G3452 (W2055, W3452);
not G3453 (W2056, W3453);
not G3454 (W2057, W3454);
not G3455 (W2058, W3455);
not G3456 (W2059, W3456);
not G3457 (W2060, W3457);
not G3458 (W2061, W3458);
not G3459 (W2062, W3459);
not G3460 (W2063, W3460);
not G3461 (W2064, W3461);
not G3462 (W2065, W3462);
not G3463 (W2066, W3463);
not G3464 (W2067, W3464);
not G3465 (W2068, W3465);
not G3466 (W2069, W3466);
not G3467 (W2070, W3467);
not G3468 (W2071, W3468);
not G3469 (W2072, W3469);
not G3470 (W2073, W3470);
not G3471 (W2074, W3471);
not G3472 (W2075, W3472);
not G3473 (W2076, W3473);
not G3474 (W2077, W3474);
not G3475 (W2078, W3475);
not G3476 (W2079, W3476);
not G3477 (W2080, W3477);
not G3478 (W2081, W3478);
not G3479 (W2082, W3479);
not G3480 (W2083, W3480);
not G3481 (W2084, W3481);
not G3482 (W2085, W3482);
not G3483 (W2086, W3483);
not G3484 (W2087, W3484);
not G3485 (W2088, W3485);
not G3486 (W2089, W3486);
not G3487 (W2090, W3487);
not G3488 (W2091, W3488);
not G3489 (W2092, W3489);
not G3490 (W2093, W3490);
not G3491 (W2094, W3491);
not G3492 (W2095, W3492);
not G3493 (W2096, W3493);
not G3494 (W2097, W3494);
not G3495 (W2098, W3495);
not G3496 (W2099, W3496);
not G3497 (W2100, W3497);
not G3498 (W2101, W3498);
not G3499 (W2102, W3499);
not G3500 (W2103, W3500);
not G3501 (W2104, W3501);
not G3502 (W2105, W3502);
not G3503 (W2106, W3503);
not G3504 (W2107, W3504);
not G3505 (W2108, W3505);
not G3506 (W2109, W3506);
not G3507 (W2110, W3507);
not G3508 (W2111, W3508);
not G3509 (W2112, W3509);
not G3510 (W2113, W3510);
not G3511 (W2114, W3511);
not G3512 (W2115, W3512);
not G3513 (W2116, W3513);
not G3514 (W2117, W3514);
not G3515 (W2118, W3515);
not G3516 (W2119, W3516);
not G3517 (W2120, W3517);
not G3518 (W2121, W3518);
not G3519 (W2122, W3519);
not G3520 (W2123, W3520);
not G3521 (W2124, W3521);
not G3522 (W2125, W3522);
not G3523 (W2126, W3523);
not G3524 (W2127, W3524);
not G3525 (W2128, W3525);
not G3526 (W2129, W3526);
not G3527 (W2130, W3527);
not G3528 (W2131, W3528);
not G3529 (W2132, W3529);
not G3530 (W2133, W3530);
not G3531 (W2134, W3531);
not G3532 (W2135, W3532);
not G3533 (W2136, W3533);
not G3534 (W2137, W3534);
not G3535 (W2138, W3535);
not G3536 (W2139, W3536);
not G3537 (W2140, W3537);
not G3538 (W2141, W3538);
not G3539 (W2142, W3539);
not G3540 (W2143, W3540);
not G3541 (W2144, W3541);
not G3542 (W2145, W3542);
not G3543 (W2146, W3543);
not G3544 (W2147, W3544);
not G3545 (W2148, W3545);
not G3546 (W2149, W3546);
not G3547 (W2150, W3547);
not G3548 (W2151, W3548);
not G3549 (W2152, W3549);
not G3550 (W2153, W3550);
not G3551 (W2154, W3551);
not G3552 (W2155, W3552);
not G3553 (W2156, W3553);
not G3554 (W2157, W3554);
not G3555 (W2158, W3555);
not G3556 (W2159, W3556);
not G3557 (W2160, W3557);
not G3558 (W2161, W3558);
not G3559 (W2162, W3559);
not G3560 (W2163, W3560);
not G3561 (W2164, W3561);
not G3562 (W2165, W3562);
not G3563 (W2166, W3563);
not G3564 (W2167, W3564);
not G3565 (W2168, W3565);
not G3566 (W2169, W3566);
not G3567 (W2170, W3567);
not G3568 (W2171, W3568);
not G3569 (W2172, W3569);
not G3570 (W2173, W3570);
not G3571 (W2174, W3571);
not G3572 (W2175, W3572);
not G3573 (W2176, W3573);
not G3574 (W2177, W3574);
not G3575 (W2178, W3575);
not G3576 (W2179, W3576);
not G3577 (W2180, W3577);
not G3578 (W2181, W3578);
not G3579 (W2182, W3579);
not G3580 (W2183, W3580);
not G3581 (W2184, W3581);
not G3582 (W2185, W3582);
not G3583 (W2186, W3583);
not G3584 (W2187, W3584);
not G3585 (W2188, W3585);
not G3586 (W2189, W3586);
not G3587 (W2190, W3587);
not G3588 (W2191, W3588);
not G3589 (W2192, W3589);
not G3590 (W2193, W3590);
not G3591 (W2194, W3591);
not G3592 (W2195, W3592);
not G3593 (W2196, W3593);
not G3594 (W2197, W3594);
not G3595 (W2198, W3595);
not G3596 (W2199, W3596);
not G3597 (W2200, W3597);
not G3598 (W2201, W3598);
not G3599 (W2202, W3599);
not G3600 (W2203, W3600);
not G3601 (W2204, W3601);
not G3602 (W2205, W3602);
not G3603 (W2206, W3603);
not G3604 (W2207, W3604);
not G3605 (W2208, W3605);
not G3606 (W2209, W3606);
not G3607 (W2210, W3607);
not G3608 (W2211, W3608);
not G3609 (W2212, W3609);
not G3610 (W2213, W3610);
not G3611 (W2214, W3611);
not G3612 (W2215, W3612);
not G3613 (W2216, W3613);
not G3614 (W2217, W3614);
not G3615 (W2218, W3615);
not G3616 (W2219, W3616);
not G3617 (W2220, W3617);
not G3618 (W2221, W3618);
not G3619 (W2222, W3619);
not G3620 (W2223, W3620);
not G3621 (W2224, W3621);
not G3622 (W2225, W3622);
not G3623 (W2226, W3623);
not G3624 (W2227, W3624);
not G3625 (W2228, W3625);
not G3626 (W2229, W3626);
not G3627 (W2230, W3627);
not G3628 (W2231, W3628);
not G3629 (W2232, W3629);
not G3630 (W2233, W3630);
not G3631 (W2234, W3631);
not G3632 (W2235, W3632);
not G3633 (W2236, W3633);
not G3634 (W2237, W3634);
not G3635 (W2238, W3635);
not G3636 (W2239, W3636);
not G3637 (W2240, W3637);
not G3638 (W2241, W3638);
not G3639 (W2242, W3639);
not G3640 (W2243, W3640);
not G3641 (W2244, W3641);
not G3642 (W2245, W3642);
not G3643 (W2246, W3643);
not G3644 (W2247, W3644);
not G3645 (W2248, W3645);
not G3646 (W2249, W3646);
not G3647 (W2250, W3647);
not G3648 (W2251, W3648);
not G3649 (W2252, W3649);
not G3650 (W2253, W3650);
not G3651 (W2254, W3651);
not G3652 (W2255, W3652);
not G3653 (W2256, W3653);
not G3654 (W2257, W3654);
not G3655 (W2258, W3655);
not G3656 (W2259, W3656);
not G3657 (W2260, W3657);
not G3658 (W2261, W3658);
not G3659 (W2262, W3659);
not G3660 (W2263, W3660);
not G3661 (W2264, W3661);
not G3662 (W2265, W3662);
not G3663 (W2266, W3663);
not G3664 (W2267, W3664);
not G3665 (W2268, W3665);
not G3666 (W2269, W3666);
not G3667 (W2270, W3667);
not G3668 (W2271, W3668);
not G3669 (W2272, W3669);
not G3670 (W2273, W3670);
not G3671 (W2274, W3671);
not G3672 (W2275, W3672);
not G3673 (W2276, W3673);
not G3674 (W2277, W3674);
not G3675 (W2278, W3675);
not G3676 (W2279, W3676);
not G3677 (W2280, W3677);
not G3678 (W2281, W3678);
not G3679 (W2282, W3679);
not G3680 (W2283, W3680);
not G3681 (W2284, W3681);
not G3682 (W2285, W3682);
not G3683 (W2286, W3683);
not G3684 (W2287, W3684);
not G3685 (W2288, W3685);
not G3686 (W2289, W3686);
not G3687 (W2290, W3687);
not G3688 (W2291, W3688);
not G3689 (W2292, W3689);
not G3690 (W2293, W3690);
not G3691 (W2294, W3691);
not G3692 (W2295, W3692);
not G3693 (W2296, W3693);
not G3694 (W2297, W3694);
not G3695 (W2298, W3695);
not G3696 (W2299, W3696);
not G3697 (W2300, W3697);
not G3698 (W2301, W3698);
not G3699 (W2302, W3699);
not G3700 (W2303, W3700);
not G3701 (W2304, W3701);
not G3702 (W2305, W3702);
not G3703 (W2306, W3703);
not G3704 (W2307, W3704);
not G3705 (W2308, W3705);
not G3706 (W2309, W3706);
not G3707 (W2310, W3707);
not G3708 (W2311, W3708);
not G3709 (W2312, W3709);
not G3710 (W2313, W3710);
not G3711 (W2314, W3711);
not G3712 (W2315, W3712);
not G3713 (W2316, W3713);
not G3714 (W2317, W3714);
not G3715 (W2318, W3715);
not G3716 (W2319, W3716);
not G3717 (W2320, W3717);
not G3718 (W2321, W3718);
not G3719 (W2322, W3719);
not G3720 (W2323, W3720);
not G3721 (W2324, W3721);
not G3722 (W2325, W3722);
not G3723 (W2326, W3723);
not G3724 (W2327, W3724);
not G3725 (W2328, W3725);
not G3726 (W2329, W3726);
not G3727 (W2330, W3727);
not G3728 (W2331, W3728);
not G3729 (W2332, W3729);
not G3730 (W2333, W3730);
not G3731 (W2334, W3731);
not G3732 (W2335, W3732);
not G3733 (W2336, W3733);
not G3734 (W2337, W3734);
not G3735 (W2338, W3735);
not G3736 (W2339, W3736);
not G3737 (W2340, W3737);
not G3738 (W2341, W3738);
not G3739 (W2342, W3739);
not G3740 (W2343, W3740);
not G3741 (W2344, W3741);
not G3742 (W2345, W3742);
not G3743 (W2346, W3743);
not G3744 (W2347, W3744);
not G3745 (W2348, W3745);
not G3746 (W2349, W3746);
not G3747 (W2350, W3747);
not G3748 (W2351, W3748);
not G3749 (W2352, W3749);
not G3750 (W2353, W3750);
not G3751 (W2354, W3751);
not G3752 (W2355, W3752);
not G3753 (W2356, W3753);
not G3754 (W2357, W3754);
not G3755 (W2358, W3755);
not G3756 (W2359, W3756);
not G3757 (W2360, W3757);
not G3758 (W2361, W3758);
not G3759 (W2362, W3759);
not G3760 (W2363, W3760);
not G3761 (W2364, W3761);
not G3762 (W2365, W3762);
not G3763 (W2366, W3763);
not G3764 (W2367, W3764);
not G3765 (W2368, W3765);
not G3766 (W2369, W3766);
not G3767 (W2370, W3767);
not G3768 (W2371, W3768);
not G3769 (W2372, W3769);
not G3770 (W2373, W3770);
not G3771 (W2374, W3771);
not G3772 (W2375, W3772);
not G3773 (W2376, W3773);
not G3774 (W2377, W3774);
not G3775 (W2378, W3775);
not G3776 (W2379, W3776);
not G3777 (W2380, W3777);
not G3778 (W2381, W3778);
not G3779 (W2382, W3779);
not G3780 (W2383, W3780);
not G3781 (W2384, W3781);
not G3782 (W2385, W3782);
not G3783 (W2386, W3783);
not G3784 (W2387, W3784);
not G3785 (W2388, W3785);
not G3786 (W2389, W3786);
not G3787 (W2390, W3787);
not G3788 (W2391, W3788);
not G3789 (W2392, W3789);
not G3790 (W2393, W3790);
not G3791 (W2394, W3791);
not G3792 (W2395, W3792);
not G3793 (W2396, W3793);
not G3794 (W2397, W3794);
not G3795 (W2398, W3795);
not G3796 (W2399, W3796);
not G3797 (W2400, W3797);
not G3798 (W2401, W3798);
not G3799 (W2402, W3799);
not G3800 (W2403, W3800);
not G3801 (W2404, W3801);
not G3802 (W2405, W3802);
not G3803 (W2406, W3803);
not G3804 (W2407, W3804);
not G3805 (W2408, W3805);
not G3806 (W2409, W3806);
not G3807 (W2410, W3807);
not G3808 (W2411, W3808);
not G3809 (W2412, W3809);
not G3810 (W2413, W3810);
not G3811 (W2414, W3811);
not G3812 (W2415, W3812);
not G3813 (W2416, W3813);
not G3814 (W2417, W3814);
not G3815 (W2418, W3815);
not G3816 (W2419, W3816);
not G3817 (W2420, W3817);
not G3818 (W2421, W3818);
not G3819 (W2422, W3819);
not G3820 (W2423, W3820);
not G3821 (W2424, W3821);
not G3822 (W2425, W3822);
not G3823 (W2426, W3823);
not G3824 (W2427, W3824);
not G3825 (W2428, W3825);
not G3826 (W2429, W3826);
not G3827 (W2430, W3827);
not G3828 (W2431, W3828);
not G3829 (W2432, W3829);
not G3830 (W2433, W3830);
not G3831 (W2434, W3831);
not G3832 (W2435, W3832);
not G3833 (W2436, W3833);
not G3834 (W2437, W3834);
not G3835 (W2438, W3835);
not G3836 (W2439, W3836);
not G3837 (W2440, W3837);
not G3838 (W2441, W3838);
not G3839 (W2442, W3839);
not G3840 (W2443, W3840);
not G3841 (W2444, W3841);
not G3842 (W2445, W3842);
not G3843 (W2446, W3843);
not G3844 (W2447, W3844);
not G3845 (W2448, W3845);
not G3846 (W2449, W3846);
not G3847 (W2450, W3847);
not G3848 (W2451, W3848);
not G3849 (W2452, W3849);
not G3850 (W2453, W3850);
not G3851 (W2454, W3851);
not G3852 (W2455, W3852);
not G3853 (W2456, W3853);
not G3854 (W2457, W3854);
not G3855 (W2458, W3855);
not G3856 (W2459, W3856);
not G3857 (W2460, W3857);
not G3858 (W2461, W3858);
not G3859 (W2462, W3859);
not G3860 (W2463, W3860);
not G3861 (W2464, W3861);
not G3862 (W2465, W3862);
not G3863 (W2466, W3863);
not G3864 (W2467, W3864);
not G3865 (W2468, W3865);
not G3866 (W2469, W3866);
not G3867 (W2470, W3867);
not G3868 (W2471, W3868);
not G3869 (W2472, W3869);
not G3870 (W2473, W3870);
not G3871 (W2474, W3871);
not G3872 (W2475, W3872);
not G3873 (W2476, W3873);
not G3874 (W2477, W3874);
not G3875 (W2478, W3875);
not G3876 (W2479, W3876);
not G3877 (W2480, W3877);
not G3878 (W2481, W3878);
not G3879 (W2482, W3879);
not G3880 (W2483, W3880);
not G3881 (W2484, W3881);
not G3882 (W2485, W3882);
not G3883 (W2486, W3883);
not G3884 (W2487, W3884);
not G3885 (W2488, W3885);
not G3886 (W2489, W3886);
not G3887 (W2490, W3887);
not G3888 (W2491, W3888);
not G3889 (W2492, W3889);
not G3890 (W2493, W3890);
not G3891 (W2494, W3891);
not G3892 (W2495, W3892);
not G3893 (W2496, W3893);
not G3894 (W2497, W3894);
not G3895 (W2498, W3895);
not G3896 (W2499, W3896);
not G3897 (W2500, W3897);
not G3898 (W2501, W3898);
not G3899 (W2502, W3899);
not G3900 (W2503, W3900);
not G3901 (W2504, W3901);
not G3902 (W2505, W3902);
not G3903 (W2506, W3903);
not G3904 (W2507, W3904);
not G3905 (W2508, W3905);
not G3906 (W2509, W3906);
not G3907 (W2510, W3907);
not G3908 (W2511, W3908);
not G3909 (W2512, W3909);
not G3910 (W2513, W3910);
not G3911 (W2514, W3911);
not G3912 (W2515, W3912);
not G3913 (W2516, W3913);
not G3914 (W2517, W3914);
not G3915 (W2518, W3915);
not G3916 (W2519, W3916);
not G3917 (W2520, W3917);
not G3918 (W2521, W3918);
not G3919 (W2522, W3919);
not G3920 (W2523, W3920);
not G3921 (W2524, W3921);
not G3922 (W2525, W3922);
not G3923 (W2526, W3923);
not G3924 (W2527, W3924);
not G3925 (W2528, W3925);
not G3926 (W2529, W3926);
not G3927 (W2530, W3927);
not G3928 (W2531, W3928);
not G3929 (W2532, W3929);
not G3930 (W2533, W3930);
not G3931 (W2534, W3931);
not G3932 (W2535, W3932);
not G3933 (W2536, W3933);
not G3934 (W2537, W3934);
not G3935 (W2538, W3935);
not G3936 (W2539, W3936);
not G3937 (W2540, W3937);
not G3938 (W2541, W3938);
not G3939 (W2542, W3939);
not G3940 (W2543, W3940);
not G3941 (W2544, W3941);
not G3942 (W2545, W3942);
not G3943 (W2546, W3943);
not G3944 (W2547, W3944);
not G3945 (W2548, W3945);
not G3946 (W2549, W3946);
not G3947 (W2550, W3947);
not G3948 (W2551, W3948);
not G3949 (W2552, W3949);
not G3950 (W2553, W3950);
not G3951 (W2554, W3951);
not G3952 (W2555, W3952);
not G3953 (W2556, W3953);
not G3954 (W2557, W3954);
not G3955 (W2558, W3955);
not G3956 (W2559, W3956);
not G3957 (W2560, W3957);
not G3958 (W2561, W3958);
not G3959 (W2562, W3959);
not G3960 (W2563, W3960);
not G3961 (W2564, W3961);
not G3962 (W2565, W3962);
not G3963 (W2566, W3963);
not G3964 (W2567, W3964);
not G3965 (W2568, W3965);
not G3966 (W2569, W3966);
not G3967 (W2570, W3967);
not G3968 (W2571, W3968);
not G3969 (W2572, W3969);
not G3970 (W2573, W3970);
not G3971 (W2574, W3971);
not G3972 (W2575, W3972);
not G3973 (W2576, W3973);
not G3974 (W2577, W3974);
not G3975 (W2578, W3975);
not G3976 (W2579, W3976);
not G3977 (W2580, W3977);
not G3978 (W2581, W3978);
not G3979 (W2582, W3979);
not G3980 (W2583, W3980);
not G3981 (W2584, W3981);
not G3982 (W2585, W3982);
not G3983 (W2586, W3983);
not G3984 (W2587, W3984);
not G3985 (W2588, W3985);
not G3986 (W2589, W3986);
not G3987 (W2590, W3987);
not G3988 (W2591, W3988);
not G3989 (W2592, W3989);
not G3990 (W2593, W3990);
not G3991 (W2594, W3991);
not G3992 (W2595, W3992);
not G3993 (W2596, W3993);
not G3994 (W2597, W3994);
not G3995 (W2598, W3995);
not G3996 (W2599, W3996);
not G3997 (W2600, W3997);
not G3998 (W2601, W3998);
not G3999 (W2602, W3999);
not G4000 (W2603, W4000);
not G4001 (W2604, W4001);
not G4002 (W2605, W4002);
not G4003 (W2606, W4003);
not G4004 (W2607, W4004);
not G4005 (W2608, W4005);
not G4006 (W2609, W4006);
not G4007 (W2610, W4007);
not G4008 (W2611, W4008);
not G4009 (W2612, W4009);
not G4010 (W2613, W4010);
not G4011 (W2614, W4011);
not G4012 (W2615, W4012);
not G4013 (W2616, W4013);
not G4014 (W2617, W4014);
not G4015 (W2618, W4015);
not G4016 (W2619, W4016);
not G4017 (W2620, W4017);
not G4018 (W2621, W4018);
not G4019 (W2622, W4019);
not G4020 (W2623, W4020);
not G4021 (W2624, W4021);
not G4022 (W2625, W4022);
not G4023 (W2626, W4023);
not G4024 (W2627, W4024);
not G4025 (W2628, W4025);
not G4026 (W2629, W4026);
not G4027 (W2630, W4027);
not G4028 (W2631, W4028);
not G4029 (W2632, W4029);
not G4030 (W2633, W4030);
not G4031 (W2634, W4031);
not G4032 (W2635, W4032);
not G4033 (W2636, W4033);
not G4034 (W2637, W4034);
not G4035 (W2638, W4035);
not G4036 (W2639, W4036);
not G4037 (W2640, W4037);
not G4038 (W2641, W4038);
not G4039 (W2642, W4039);
not G4040 (W2643, W4040);
not G4041 (W2644, W4041);
not G4042 (W2645, W4042);
not G4043 (W2646, W4043);
not G4044 (W2647, W4044);
not G4045 (W2648, W4045);
not G4046 (W2649, W4046);
not G4047 (W2650, W4047);
not G4048 (W2651, W4048);
not G4049 (W2652, W4049);
not G4050 (W2653, W4050);
not G4051 (W2654, W4051);
not G4052 (W2655, W4052);
not G4053 (W2656, W4053);
not G4054 (W2657, W4054);
not G4055 (W2658, W4055);
not G4056 (W2659, W4056);
not G4057 (W2660, W4057);
not G4058 (W2661, W4058);
not G4059 (W2662, W4059);
not G4060 (W2663, W4060);
not G4061 (W2664, W4061);
not G4062 (W2665, W4062);
not G4063 (W2666, W4063);
not G4064 (W2667, W4064);
not G4065 (W2668, W4065);
not G4066 (W2669, W4066);
not G4067 (W2670, W4067);
not G4068 (W2671, W4068);
not G4069 (W2672, W4069);
not G4070 (W2673, W4070);
not G4071 (W2674, W4071);
not G4072 (W2675, W4072);
not G4073 (W2676, W4073);
not G4074 (W2677, W4074);
not G4075 (W2678, W4075);
not G4076 (W2679, W4076);
not G4077 (W2680, W4077);
not G4078 (W2681, W4078);
not G4079 (W2682, W4079);
not G4080 (W2683, W4080);
not G4081 (W2684, W4081);
not G4082 (W2685, W4082);
not G4083 (W2686, W4083);
not G4084 (W2687, W4084);
not G4085 (W2688, W4085);
not G4086 (W2689, W4086);
not G4087 (W2690, W4087);
not G4088 (W2691, W4088);
not G4089 (W2692, W4089);
not G4090 (W2693, W4090);
not G4091 (W2694, W4091);
not G4092 (W2695, W4092);
not G4093 (W2696, W4093);
not G4094 (W2697, W4094);
not G4095 (W2698, W4095);
not G4096 (W2699, W4096);
not G4097 (W2700, W4097);
not G4098 (W2701, W4098);
not G4099 (W2702, W4099);
not G4100 (W2703, W4100);
not G4101 (W2704, W4101);
not G4102 (W2705, W4102);
not G4103 (W2706, W4103);
not G4104 (W2707, W4104);
not G4105 (W2708, W4105);
not G4106 (W2709, W4106);
not G4107 (W2710, W4107);
not G4108 (W2711, W4108);
not G4109 (W2712, W4109);
not G4110 (W2713, W4110);
not G4111 (W2714, W4111);
not G4112 (W2715, W4112);
not G4113 (W2716, W4113);
not G4114 (W2717, W4114);
not G4115 (W2718, W4115);
not G4116 (W2719, W4116);
not G4117 (W2720, W4117);
not G4118 (W2721, W4118);
not G4119 (W2722, W4119);
not G4120 (W2723, W4120);
not G4121 (W2724, W4121);
not G4122 (W2725, W4122);
not G4123 (W2726, W4123);
not G4124 (W2727, W4124);
not G4125 (W2728, W4125);
not G4126 (W2729, W4126);
not G4127 (W2730, W4127);
not G4128 (W2731, W4128);
not G4129 (W2732, W4129);
not G4130 (W2733, W4130);
not G4131 (W2734, W4131);
not G4132 (W2735, W4132);
not G4133 (W2736, W4133);
not G4134 (W2737, W4134);
not G4135 (W2738, W4135);
not G4136 (W2739, W4136);
not G4137 (W2740, W4137);
not G4138 (W2741, W4138);
not G4139 (W2742, W4139);
not G4140 (W2743, W4140);
not G4141 (W2744, W4141);
not G4142 (W2745, W4142);
not G4143 (W2746, W4143);
not G4144 (W2747, W4144);
not G4145 (W2748, W4145);
not G4146 (W2749, W4146);
not G4147 (W2750, W4147);
not G4148 (W2751, W4148);
not G4149 (W2752, W4149);
not G4150 (W2753, W4150);
not G4151 (W2754, W4151);
not G4152 (W2755, W4152);
not G4153 (W2756, W4153);
not G4154 (W2757, W4154);
not G4155 (W2758, W4155);
not G4156 (W2759, W4156);
not G4157 (W2760, W4157);
not G4158 (W2761, W4158);
not G4159 (W2762, W4159);
not G4160 (W2763, W4160);
not G4161 (W2764, W4161);
not G4162 (W2765, W4162);
not G4163 (W2766, W4163);
not G4164 (W2767, W4164);
not G4165 (W2768, W4165);
not G4166 (W2769, W4166);
not G4167 (W2770, W4167);
not G4168 (W2771, W4168);
not G4169 (W2772, W4169);
not G4170 (W2773, W4170);
not G4171 (W2774, W4171);
not G4172 (W2775, W4172);
not G4173 (W2776, W4173);
not G4174 (W2777, W4174);
not G4175 (W2778, W4175);
not G4176 (W2779, W4176);
not G4177 (W2780, W4177);
not G4178 (W2781, W4178);
not G4179 (W2782, W4179);
not G4180 (W2783, W4180);
not G4181 (W2784, W4181);
not G4182 (W2785, W4182);
not G4183 (W2786, W4183);
not G4184 (W2787, W4184);
not G4185 (W2788, W4185);
not G4186 (W2789, W4186);
not G4187 (W2790, W4187);
not G4188 (W2791, W4188);
not G4189 (W2792, W4189);
not G4190 (W2793, W4190);
not G4191 (W2794, W4191);
not G4192 (W2795, W4192);
not G4193 (W2796, W4192);
not G4194 (W2797, W4192);
not G4195 (W2798, W4192);
not G4196 (W2799, W4193);
not G4197 (W2800, W4194);
not G4198 (W2801, W4194);
not G4199 (W2802, W4194);
not G4200 (W2803, W4195);
not G4201 (W2804, W4196);
not G4202 (W2805, W4197);
not G4203 (W2806, W4198);
not G4204 (W2807, W4199);
not G4205 (W2808, W4200);
not G4206 (W2809, W4201);
not G4207 (W2810, W4202);
not G4208 (W2811, W4203);
not G4209 (W2812, W4204);
not G4210 (W2813, W4205);
not G4211 (W2814, W4206);
not G4212 (W2815, W4207);
not G4213 (W2816, W4208);
not G4214 (W2817, W4209);
not G4215 (W2818, W4210);
not G4216 (W2819, W4211);
not G4217 (W2820, W4212);
not G4218 (W2821, W4213);
not G4219 (W2822, W4214);
not G4220 (W2823, W4215);
not G4221 (W2824, W4216);
not G4222 (W2825, W4217);
not G4223 (W2826, W4218);
not G4224 (W2827, W4219);
not G4225 (W2828, W4220);
not G4226 (W2829, W4221);
not G4227 (W2830, W4222);
not G4228 (W2831, W4223);
not G4229 (W2832, W4224);
not G4230 (W2833, W4225);
not G4231 (W2834, W4226);
not G4232 (W2835, W4227);
not G4233 (W2836, W4228);
not G4234 (W2837, W4229);
not G4235 (W2838, W4230);
not G4236 (W2839, W4231);
not G4237 (W2840, W4232);
not G4238 (W2841, W4233);
not G4239 (W2842, W4234);
not G4240 (W2843, W4235);
not G4241 (W2844, W4236);
not G4242 (W2845, W4237);
not G4243 (W2846, W4238);
not G4244 (W2847, W4239);
not G4245 (W2848, W4240);
not G4246 (W2849, W4241);
not G4247 (W2850, W4242);
not G4248 (W2851, W4243);
not G4249 (W2852, W4244);
not G4250 (W2853, W4245);
not G4251 (W2854, W4246);
not G4252 (W2855, W4247);
not G4253 (W2856, W4248);
not G4254 (W2857, W4249);
not G4255 (W2858, W4250);
not G4256 (W2859, W4251);
not G4257 (W2860, W4252);
not G4258 (W2861, W4253);
not G4259 (W2862, W4254);
not G4260 (W2863, W4255);
not G4261 (W2864, W4256);
not G4262 (W2865, W4257);
not G4263 (W2866, W4258);
not G4264 (W2867, W4259);
not G4265 (W2868, W4260);
not G4266 (W2869, W4261);
not G4267 (W2870, W4262);
not G4268 (W2871, W4263);
not G4269 (W2872, W4264);
not G4270 (W2873, W4265);
not G4271 (W2874, W4266);
not G4272 (W2875, W4267);
not G4273 (W2876, W4268);
not G4274 (W2877, W4269);
not G4275 (W2878, W4270);
not G4276 (W2879, W4271);
not G4277 (W2880, W4272);
not G4278 (W2881, W4273);
not G4279 (W2882, W4274);
not G4280 (W2883, W4275);
not G4281 (W2884, W4276);
not G4282 (W2885, W4277);
not G4283 (W2886, W4278);
not G4284 (W2887, W4279);
not G4285 (W2888, W4280);
not G4286 (W2889, W4281);
not G4287 (W2890, W4282);
not G4288 (W2891, W4283);
not G4289 (W2892, W4284);
not G4290 (W2893, W4285);
not G4291 (W2894, W4286);
not G4292 (W2895, W4287);
not G4293 (W2896, W4288);
not G4294 (W2897, W4289);
not G4295 (W2898, W4290);
not G4296 (W2899, W4291);
not G4297 (W2900, W4292);
not G4298 (W2901, W4293);
not G4299 (W2902, W4294);
not G4300 (W2903, W4295);
not G4301 (W2904, W4296);
not G4302 (W2905, W4297);
not G4303 (W2906, W4298);
not G4304 (W2907, W4299);
not G4305 (W2908, W4300);
not G4306 (W2909, W4301);
not G4307 (W2910, W4302);
not G4308 (W2911, W4303);
not G4309 (W2912, W4304);
not G4310 (W2913, W4305);
not G4311 (W2914, W4306);
not G4312 (W2915, W4307);
not G4313 (W2916, W4308);
not G4314 (W2917, W4309);
not G4315 (W2918, W4310);
not G4316 (W2919, W4311);
not G4317 (W2920, W4312);
not G4318 (W2921, W4313);
not G4319 (W2922, W4314);
not G4320 (W2923, W4315);
not G4321 (W2924, W4316);
not G4322 (W2925, W4317);
not G4323 (W2926, W4318);
not G4324 (W2927, W4319);
not G4325 (W2928, W4320);
not G4326 (W2929, W4321);
not G4327 (W2930, W4322);
not G4328 (W2931, W4323);
not G4329 (W2932, W4324);
not G4330 (W2933, W4325);
not G4331 (W2934, W4326);
not G4332 (W2935, W4327);
not G4333 (W2936, W4328);
not G4334 (W2937, W4329);
not G4335 (W2938, W4330);
not G4336 (W2939, W4331);
not G4337 (W2940, W4332);
not G4338 (W2941, W4333);
not G4339 (W2942, W4334);
not G4340 (W2943, W4335);
not G4341 (W2944, W4336);
not G4342 (W2945, W4337);
not G4343 (W2946, W4338);
not G4344 (W2947, W4339);
not G4345 (W2948, W4340);
not G4346 (W2949, W4341);
not G4347 (W2950, W4342);
not G4348 (W2951, W4343);
not G4349 (W2952, W4344);
not G4350 (W2953, W4345);
not G4351 (W2954, W4346);
not G4352 (W2955, W4347);
not G4353 (W2956, W4348);
not G4354 (W2957, W4349);
not G4355 (W2958, W4350);
not G4356 (W2959, W4351);
not G4357 (W2960, W4352);
not G4358 (W2961, W4353);
not G4359 (W2962, W4354);
not G4360 (W2963, W4355);
not G4361 (W2964, W4356);
not G4362 (W2965, W4357);
not G4363 (W2966, W4358);
not G4364 (W2967, W4359);
not G4365 (W2968, W4360);
not G4366 (W2969, W4361);
not G4367 (W2970, W4362);
not G4368 (W2971, W4363);
not G4369 (W2972, W4364);
not G4370 (W2973, W4365);
not G4371 (W2974, W4366);
not G4372 (W2975, W4367);
not G4373 (W2976, W4368);
not G4374 (W2977, W4369);
not G4375 (W2978, W4370);
not G4376 (W2979, W4371);
not G4377 (W2980, W4372);
not G4378 (W2981, W4373);
not G4379 (W2982, W4374);
not G4380 (W2983, W4375);
not G4381 (W2984, W4376);
not G4382 (W2985, W4377);
not G4383 (W2986, W4378);
not G4384 (W2987, W4379);
not G4385 (W2988, W4380);
not G4386 (W2989, W4381);
not G4387 (W2990, W4382);
not G4388 (W2991, W4383);
not G4389 (W2992, W4384);
not G4390 (W2993, W4385);
not G4391 (W2994, W4386);
not G4392 (W2995, W4387);
not G4393 (W2996, W4388);
not G4394 (W2997, W4389);
not G4395 (W2998, W4390);
not G4396 (W2999, W4391);
not G4397 (W3000, W4392);
not G4398 (W3001, W4393);
not G4399 (W3002, W4394);
not G4400 (W3003, W4395);
not G4401 (W3004, W4396);
not G4402 (W3005, W4397);
not G4403 (W3006, W4398);
not G4404 (W3007, W4399);
not G4405 (W3008, W4400);
not G4406 (W3009, W4401);
not G4407 (W3010, W4402);
not G4408 (W3011, W4403);
not G4409 (W3012, W4404);
not G4410 (W3013, W4405);
not G4411 (W3014, W4406);
not G4412 (W3015, W4407);
not G4413 (W3016, W4408);
not G4414 (W3017, W4409);
not G4415 (W3018, W4410);
not G4416 (W3019, W4411);
not G4417 (W3020, W4412);
not G4418 (W3021, W4413);
not G4419 (W3022, W4414);
not G4420 (W3023, W4415);
not G4421 (W3024, W4416);
not G4422 (W3025, W4417);
not G4423 (W3026, W4418);
not G4424 (W3027, W4419);
not G4425 (W3028, W4420);
not G4426 (W3029, W4421);
not G4427 (W3030, W4422);
not G4428 (W3031, W4423);
not G4429 (W3032, W4424);
not G4430 (W3033, W4425);
not G4431 (W3034, W4426);
not G4432 (W3035, W4427);
not G4433 (W3036, W4428);
not G4434 (W3037, W4429);
not G4435 (W3038, W4430);
not G4436 (W3039, W4431);
not G4437 (W3040, W4432);
not G4438 (W3041, W4433);
not G4439 (W3042, W4434);
not G4440 (W3043, W4435);
not G4441 (W3044, W4436);
not G4442 (W3045, W4437);
not G4443 (W3046, W4438);
not G4444 (W3047, I219);
not G4445 (W3048, W4439);
not G4446 (W3049, W4440);
not G4447 (W3050, W4441);
not G4448 (W3051, W4442);
not G4449 (W3052, W4443);
not G4450 (W3053, W4444);
not G4451 (W3054, W4445);
not G4452 (W3055, W4446);
not G4453 (W3056, W4447);
not G4454 (W3057, W4448);
not G4455 (W3058, W4449);
not G4456 (W3059, W4450);
not G4457 (W3060, W4451);
not G4458 (W3061, W4452);
not G4459 (W3062, W4453);
not G4460 (W3063, W4454);
not G4461 (W3064, W4455);
not G4462 (W3065, W4456);
not G4463 (W3066, W4457);
not G4464 (W3067, W4458);
not G4465 (W3068, W4459);
not G4466 (W3069, W4460);
not G4467 (W3070, W4461);
not G4468 (W3071, W4462);
not G4469 (W3072, W4463);
not G4470 (W3073, W4464);
not G4471 (W3074, W4465);
not G4472 (W3075, W4466);
not G4473 (W3076, W4467);
not G4474 (W3077, W4468);
not G4475 (W3078, W4469);
not G4476 (W3079, W4470);
not G4477 (W3080, W4471);
not G4478 (W3081, W4472);
not G4479 (W3082, W4473);
not G4480 (W3083, W4474);
not G4481 (W3084, W4475);
not G4482 (W3085, W4476);
not G4483 (W3086, W4477);
not G4484 (W3087, W4478);
not G4485 (W3088, W4479);
not G4486 (W3089, W4480);
not G4487 (W3090, W4481);
not G4488 (W3091, W4482);
not G4489 (W3092, W4483);
not G4490 (W3093, W4484);
not G4491 (W3094, W4485);
not G4492 (W3095, W4486);
not G4493 (W3096, W4487);
not G4494 (W3097, W4488);
not G4495 (W3098, W4489);
not G4496 (W3099, W4490);
not G4497 (W3100, W4491);
not G4498 (W3101, W4492);
not G4499 (W3102, W4493);
not G4500 (W3103, W4494);
not G4501 (W3104, W4495);
not G4502 (W3105, W4496);
not G4503 (W3106, W4497);
not G4504 (W3107, W4498);
not G4505 (W3108, W4499);
not G4506 (W3109, W4500);
not G4507 (W3110, W4501);
not G4508 (W3111, W4502);
not G4509 (W3112, W4503);
not G4510 (W3113, W4504);
not G4511 (W3114, W4505);
not G4512 (W3115, W4506);
not G4513 (W3116, W4507);
not G4514 (W3117, W4508);
not G4515 (W3118, W4509);
not G4516 (W3119, W4510);
not G4517 (W3120, W4511);
not G4518 (W3121, W4512);
not G4519 (W3122, W4513);
not G4520 (W3123, W4514);
not G4521 (W3124, W4515);
not G4522 (W3125, W4516);
not G4523 (W3126, W4517);
not G4524 (W3127, W4518);
not G4525 (W3128, W4519);
not G4526 (W3129, W4520);
not G4527 (W3130, W4521);
not G4528 (W3131, W4522);
not G4529 (W3132, W4523);
not G4530 (W3133, W4524);
not G4531 (W3134, W4525);
not G4532 (W3135, W4526);
not G4533 (W3136, W4527);
not G4534 (W3137, W4528);
not G4535 (W3138, W4529);
not G4536 (W3139, W4530);
not G4537 (W3140, W4531);
not G4538 (W3141, W4532);
not G4539 (W3142, W4533);
not G4540 (W3143, W4534);
not G4541 (W3144, W4535);
not G4542 (W3145, W4536);
not G4543 (W3146, W4537);
not G4544 (W3147, W4538);
not G4545 (W3148, W4539);
not G4546 (W3149, W4540);
not G4547 (W3150, W4541);
not G4548 (W3151, W4542);
not G4549 (W3152, W4543);
not G4550 (W3153, W4544);
not G4551 (W3154, W4545);
not G4552 (W3155, W4546);
not G4553 (W3156, W4547);
not G4554 (W3157, W4548);
not G4555 (W3158, W4549);
not G4556 (W3159, W4550);
not G4557 (W3160, W4551);
not G4558 (W3161, W4552);
not G4559 (W3162, W4553);
not G4560 (W3163, W4554);
not G4561 (W3164, W4555);
not G4562 (W3165, W4556);
not G4563 (W3166, W4557);
not G4564 (W3167, W4558);
not G4565 (W3168, W4559);
not G4566 (W3169, W4560);
not G4567 (W3170, W4561);
not G4568 (W3171, W4562);
not G4569 (W3172, W4563);
not G4570 (W3173, W4564);
not G4571 (W3174, W4565);
not G4572 (W3175, W4566);
not G4573 (W3176, W4567);
not G4574 (W3177, W4568);
not G4575 (W3178, W4569);
not G4576 (W3179, W4570);
not G4577 (W3180, W4571);
not G4578 (W3181, W4572);
not G4579 (W3182, W4573);
not G4580 (W3183, W4574);
not G4581 (W3184, W4575);
not G4582 (W3185, W4576);
not G4583 (W3186, W4577);
not G4584 (W3187, W4578);
not G4585 (W3188, W4579);
not G4586 (W3189, W4580);
not G4587 (W3190, W4581);
not G4588 (W3191, W4582);
not G4589 (W3192, W4583);
not G4590 (W3193, W4584);
not G4591 (W3194, W4585);
not G4592 (W3195, W4586);
not G4593 (W3196, W4587);
not G4594 (W3197, W4588);
not G4595 (W3198, W4589);
not G4596 (W3199, W4590);
not G4597 (W3200, W4591);
not G4598 (W3201, W4592);
not G4599 (W3202, W4593);
not G4600 (W3203, W4594);
not G4601 (W3204, W4595);
not G4602 (W3205, W4596);
not G4603 (W3206, W4597);
not G4604 (W3207, W4598);
not G4605 (W3208, W4599);
not G4606 (W3209, W4600);
not G4607 (W3210, W4601);
not G4608 (W3211, W4602);
not G4609 (W3212, W4603);
not G4610 (W3213, W4604);
not G4611 (W3214, W4605);
not G4612 (W3215, W4606);
not G4613 (W3216, W4607);
not G4614 (W3217, W4608);
not G4615 (W3218, W4609);
not G4616 (W3219, W4610);
not G4617 (W3220, W4611);
not G4618 (W3221, W4612);
not G4619 (W3222, W4613);
not G4620 (W3223, W4614);
not G4621 (W3224, W4615);
not G4622 (W3225, W4616);
not G4623 (W3226, W4617);
not G4624 (W3227, W4618);
not G4625 (W3228, W4619);
not G4626 (W3229, W4620);
not G4627 (W3230, W4621);
not G4628 (W3231, W4622);
not G4629 (W3232, W4623);
not G4630 (W3233, W4624);
not G4631 (W3234, W4625);
not G4632 (W3235, W4626);
not G4633 (W3236, W4627);
not G4634 (W3237, W4628);
not G4635 (W3238, W4629);
not G4636 (W3239, W4630);
not G4637 (W3240, W4631);
not G4638 (W3241, W4632);
not G4639 (W3242, W4633);
not G4640 (W3243, W4634);
not G4641 (W3244, W4635);
not G4642 (W3245, W4636);
not G4643 (W3246, W4637);
not G4644 (W3247, W4638);
not G4645 (W3248, W4639);
not G4646 (W3249, W4640);
not G4647 (W3250, W4641);
not G4648 (W3251, W4642);
not G4649 (W3252, W4643);
not G4650 (W3253, W4644);
not G4651 (W3254, W4645);
not G4652 (W3255, W4646);
not G4653 (W3256, W4647);
not G4654 (W3257, W4648);
not G4655 (W3258, W4649);
not G4656 (W3259, W4650);
not G4657 (W3260, W4651);
not G4658 (W3261, W4652);
not G4659 (W3262, W4653);
not G4660 (W3263, W4654);
not G4661 (W3264, W4655);
not G4662 (W3265, W4656);
not G4663 (W3266, W4657);
not G4664 (W3267, W4658);
not G4665 (W3268, W4659);
not G4666 (W3269, W4660);
not G4667 (W3270, W4661);
not G4668 (W3271, W4662);
not G4669 (W3272, W4663);
not G4670 (W3273, W4664);
not G4671 (W3274, W4665);
not G4672 (W3275, W4666);
not G4673 (W3276, W4667);
not G4674 (W3277, W4668);
not G4675 (W3278, W4669);
not G4676 (W3279, W4670);
not G4677 (W3280, W4671);
not G4678 (W3281, W4672);
not G4679 (W3282, W4673);
not G4680 (W3283, W4674);
not G4681 (W3284, W4675);
not G4682 (W3285, W4676);
not G4683 (W3286, W4677);
not G4684 (W3287, W4678);
not G4685 (W3288, W4679);
not G4686 (W3289, W4680);
not G4687 (W3290, W4681);
not G4688 (W3291, W4682);
not G4689 (W3292, W4683);
not G4690 (W3293, W4684);
not G4691 (W3294, W4685);
not G4692 (W3295, W4686);
not G4693 (W3296, W4687);
not G4694 (W3297, W4688);
not G4695 (W3298, W4689);
not G4696 (W3299, W4690);
not G4697 (W3300, W4691);
not G4698 (W3301, W4692);
not G4699 (W3302, W4693);
not G4700 (W3303, W4694);
not G4701 (W3304, W4695);
not G4702 (W3305, W4696);
not G4703 (W3306, W4697);
not G4704 (W3307, W4698);
not G4705 (W3308, W4699);
not G4706 (W3309, W4700);
not G4707 (W3310, W4701);
not G4708 (W3311, W4702);
not G4709 (W3312, W4703);
not G4710 (W3313, W4704);
not G4711 (W3314, W4705);
not G4712 (W3315, W4706);
not G4713 (W3316, W4707);
not G4714 (W3317, W4708);
not G4715 (W3318, W4709);
not G4716 (W3319, W4710);
not G4717 (W3320, W4711);
not G4718 (W3321, W4712);
not G4719 (W3322, W4713);
not G4720 (W3323, I220);
not G4721 (W3324, W4714);
not G4722 (W3325, W4715);
not G4723 (W3326, W4716);
not G4724 (W3327, W4717);
not G4725 (W3328, W4718);
not G4726 (W3329, W4719);
not G4727 (W3330, W4720);
not G4728 (W3331, W4721);
not G4729 (W3332, W4722);
not G4730 (W3333, W4723);
not G4731 (W3334, W4724);
not G4732 (W3335, W4725);
not G4733 (W3336, W4726);
not G4734 (W3337, W4727);
not G4735 (W3338, W4728);
not G4736 (W3339, W4729);
not G4737 (W3340, W4730);
not G4738 (W3341, W4731);
not G4739 (W3342, W4732);
not G4740 (W3343, W4733);
not G4741 (W3344, W4734);
not G4742 (W3345, W4735);
not G4743 (W3346, W4736);
not G4744 (W3347, W4737);
not G4745 (W3348, W4738);
not G4746 (W3349, W4739);
not G4747 (W3350, W4740);
not G4748 (W3351, W4741);
not G4749 (W3352, W4742);
not G4750 (W3353, W4743);
not G4751 (W3354, W4744);
not G4752 (W3355, W4745);
not G4753 (W3356, W4746);
not G4754 (W3357, W4747);
not G4755 (W3358, W4748);
not G4756 (W3359, W4749);
not G4757 (W3360, W4750);
not G4758 (W3361, W4751);
not G4759 (W3362, W4752);
not G4760 (W3363, W4753);
not G4761 (W3364, W4754);
not G4762 (W3365, W4755);
not G4763 (W3366, W4756);
not G4764 (W3367, W4757);
not G4765 (W3368, W4758);
not G4766 (W3369, W4759);
not G4767 (W3370, W4760);
not G4768 (W3371, W4761);
not G4769 (W3372, W4762);
not G4770 (W3373, W4763);
not G4771 (W3374, W4764);
not G4772 (W3375, W4765);
not G4773 (W3376, W4766);
not G4774 (W3377, W4767);
not G4775 (W3378, W4768);
not G4776 (W3379, W4769);
not G4777 (W3380, W4770);
not G4778 (W3381, W4771);
not G4779 (W3382, W4772);
not G4780 (W3383, W4773);
not G4781 (W3384, W4774);
not G4782 (W3385, W4775);
not G4783 (W3386, W4776);
not G4784 (W3387, W4777);
not G4785 (W3388, W4778);
not G4786 (W3389, W4779);
not G4787 (W3390, W4780);
not G4788 (W3391, W4781);
not G4789 (W3392, W4782);
not G4790 (W3393, W4783);
not G4791 (W3394, W4784);
not G4792 (W3395, W4785);
not G4793 (W3396, W4786);
not G4794 (W3397, W4787);
not G4795 (W3398, W4788);
not G4796 (W3399, W4789);
not G4797 (W3400, W4790);
not G4798 (W3401, W4791);
not G4799 (W3402, W4792);
not G4800 (W3403, W4793);
not G4801 (W3404, W4794);
not G4802 (W3405, W4795);
not G4803 (W3406, W4796);
not G4804 (W3407, W4797);
not G4805 (W3408, W4798);
not G4806 (W3409, W4799);
not G4807 (W3410, W4800);
not G4808 (W3411, W4801);
not G4809 (W3412, W4802);
not G4810 (W3413, W4803);
not G4811 (W3414, W4804);
not G4812 (W3415, W4805);
not G4813 (W3416, W4806);
not G4814 (W3417, W4807);
not G4815 (W3418, W4808);
not G4816 (W3419, W4809);
not G4817 (W3420, W4810);
not G4818 (W3421, W4811);
not G4819 (W3422, W4812);
not G4820 (W3423, W4813);
not G4821 (W3424, W4814);
not G4822 (W3425, W4815);
not G4823 (W3426, W4816);
not G4824 (W3427, W4817);
not G4825 (W3428, W4818);
not G4826 (W3429, W4819);
not G4827 (W3430, W4820);
not G4828 (W3431, W4821);
not G4829 (W3432, W4822);
not G4830 (W3433, W4823);
not G4831 (W3434, W4824);
not G4832 (W3435, W4825);
not G4833 (W3436, W4826);
not G4834 (W3437, W4827);
not G4835 (W3438, W4828);
not G4836 (W3439, W4829);
not G4837 (W3440, W4830);
not G4838 (W3441, W4831);
not G4839 (W3442, W4832);
not G4840 (W3443, W4833);
not G4841 (W3444, W4834);
not G4842 (W3445, W4835);
not G4843 (W3446, W4836);
not G4844 (W3447, W4837);
not G4845 (W3448, W4838);
not G4846 (W3449, W4839);
not G4847 (W3450, W4840);
not G4848 (W3451, W4841);
not G4849 (W3452, W4842);
not G4850 (W3453, W4843);
not G4851 (W3454, W4844);
not G4852 (W3455, W4845);
not G4853 (W3456, W4846);
not G4854 (W3457, W4847);
not G4855 (W3458, W4848);
not G4856 (W3459, W4849);
not G4857 (W3460, W4850);
not G4858 (W3461, W4851);
not G4859 (W3462, W4852);
not G4860 (W3463, W4853);
not G4861 (W3464, W4854);
not G4862 (W3465, W4855);
not G4863 (W3466, W4856);
not G4864 (W3467, W4857);
not G4865 (W3468, W4858);
not G4866 (W3469, W4859);
not G4867 (W3470, W4860);
not G4868 (W3471, W4861);
not G4869 (W3472, W4862);
not G4870 (W3473, W4863);
not G4871 (W3474, W4864);
not G4872 (W3475, W4865);
not G4873 (W3476, W4866);
not G4874 (W3477, W4867);
not G4875 (W3478, W4868);
not G4876 (W3479, W4869);
not G4877 (W3480, W4870);
not G4878 (W3481, W4871);
not G4879 (W3482, W4872);
not G4880 (W3483, W4873);
not G4881 (W3484, W4874);
not G4882 (W3485, W4875);
not G4883 (W3486, W4876);
not G4884 (W3487, W4877);
not G4885 (W3488, W4878);
not G4886 (W3489, W4879);
not G4887 (W3490, W4880);
not G4888 (W3491, W4881);
not G4889 (W3492, W4882);
not G4890 (W3493, W4883);
not G4891 (W3494, W4884);
not G4892 (W3495, W4885);
not G4893 (W3496, W4886);
not G4894 (W3497, W4887);
not G4895 (W3498, W4888);
not G4896 (W3499, W4889);
not G4897 (W3500, W4890);
not G4898 (W3501, W4891);
not G4899 (W3502, W4892);
not G4900 (W3503, W4893);
not G4901 (W3504, W4894);
not G4902 (W3505, W4895);
not G4903 (W3506, W4896);
not G4904 (W3507, W4897);
not G4905 (W3508, W4898);
not G4906 (W3509, W4899);
not G4907 (W3510, W4900);
not G4908 (W3511, W4901);
not G4909 (W3512, W4902);
not G4910 (W3513, W4903);
not G4911 (W3514, W4904);
not G4912 (W3515, W4905);
not G4913 (W3516, W4906);
not G4914 (W3517, W4907);
not G4915 (W3518, W4908);
not G4916 (W3519, W4909);
not G4917 (W3520, W4910);
not G4918 (W3521, W4911);
not G4919 (W3522, W4912);
not G4920 (W3523, W4913);
not G4921 (W3524, W4914);
not G4922 (W3525, W4915);
not G4923 (W3526, W4916);
not G4924 (W3527, W4917);
not G4925 (W3528, W4918);
not G4926 (W3529, W4919);
not G4927 (W3530, W4920);
not G4928 (W3531, W4921);
not G4929 (W3532, W4922);
not G4930 (W3533, W4923);
not G4931 (W3534, W4924);
not G4932 (W3535, W4925);
not G4933 (W3536, W4926);
not G4934 (W3537, W4927);
not G4935 (W3538, W4928);
not G4936 (W3539, W4929);
not G4937 (W3540, W4930);
not G4938 (W3541, W4931);
not G4939 (W3542, W4932);
not G4940 (W3543, W4933);
not G4941 (W3544, W4934);
not G4942 (W3545, W4935);
not G4943 (W3546, W4936);
not G4944 (W3547, W4937);
not G4945 (W3548, W4938);
not G4946 (W3549, W4939);
not G4947 (W3550, W4940);
not G4948 (W3551, W4941);
not G4949 (W3552, W4942);
not G4950 (W3553, W4943);
not G4951 (W3554, W4944);
not G4952 (W3555, W4945);
not G4953 (W3556, W4946);
not G4954 (W3557, W4947);
not G4955 (W3558, W4948);
not G4956 (W3559, W4949);
not G4957 (W3560, W4950);
not G4958 (W3561, W4951);
not G4959 (W3562, W4952);
not G4960 (W3563, W4953);
not G4961 (W3564, W4954);
not G4962 (W3565, W4955);
not G4963 (W3566, W4956);
not G4964 (W3567, W4957);
not G4965 (W3568, W4958);
not G4966 (W3569, W4959);
not G4967 (W3570, W4960);
not G4968 (W3571, W4961);
not G4969 (W3572, W4962);
not G4970 (W3573, W4963);
not G4971 (W3574, W4964);
not G4972 (W3575, W4965);
not G4973 (W3576, W4966);
not G4974 (W3577, W4967);
not G4975 (W3578, W4968);
not G4976 (W3579, W4969);
not G4977 (W3580, W4970);
not G4978 (W3581, W4971);
not G4979 (W3582, W4972);
not G4980 (W3583, W4973);
not G4981 (W3584, W4974);
not G4982 (W3585, W4975);
not G4983 (W3586, W4976);
not G4984 (W3587, W4977);
not G4985 (W3588, W4978);
not G4986 (W3589, W4979);
not G4987 (W3590, W4980);
not G4988 (W3591, W4981);
not G4989 (W3592, W4982);
not G4990 (W3593, W4983);
not G4991 (W3594, W4984);
not G4992 (W3595, W4985);
not G4993 (W3596, W4986);
not G4994 (W3597, W4987);
not G4995 (W3598, W4988);
not G4996 (W3599, I221);
not G4997 (W3600, W4989);
not G4998 (W3601, W4990);
not G4999 (W3602, W4991);
not G5000 (W3603, W4992);
not G5001 (W3604, W4993);
not G5002 (W3605, W4994);
not G5003 (W3606, W4995);
not G5004 (W3607, W4996);
not G5005 (W3608, W4997);
not G5006 (W3609, W4998);
not G5007 (W3610, W4999);
not G5008 (W3611, W5000);
not G5009 (W3612, W5001);
not G5010 (W3613, W5002);
not G5011 (W3614, W5003);
not G5012 (W3615, W5004);
not G5013 (W3616, W5005);
not G5014 (W3617, W5006);
not G5015 (W3618, W5007);
not G5016 (W3619, W5008);
not G5017 (W3620, W5009);
not G5018 (W3621, W5010);
not G5019 (W3622, W5011);
not G5020 (W3623, W5012);
not G5021 (W3624, W5013);
not G5022 (W3625, W5014);
not G5023 (W3626, W5015);
not G5024 (W3627, W5016);
not G5025 (W3628, W5017);
not G5026 (W3629, W5018);
not G5027 (W3630, W5019);
not G5028 (W3631, W5020);
not G5029 (W3632, W5021);
not G5030 (W3633, W5022);
not G5031 (W3634, W5023);
not G5032 (W3635, W5024);
not G5033 (W3636, W5025);
not G5034 (W3637, W5026);
not G5035 (W3638, W5027);
not G5036 (W3639, W5028);
not G5037 (W3640, W5029);
not G5038 (W3641, W5030);
not G5039 (W3642, W5031);
not G5040 (W3643, W5032);
not G5041 (W3644, W5033);
not G5042 (W3645, W5034);
not G5043 (W3646, W5035);
not G5044 (W3647, W5036);
not G5045 (W3648, W5037);
not G5046 (W3649, W5038);
not G5047 (W3650, W5039);
not G5048 (W3651, W5040);
not G5049 (W3652, W5041);
not G5050 (W3653, W5042);
not G5051 (W3654, W5043);
not G5052 (W3655, W5044);
not G5053 (W3656, W5045);
not G5054 (W3657, W5046);
not G5055 (W3658, W5047);
not G5056 (W3659, W5048);
not G5057 (W3660, W5049);
not G5058 (W3661, W5050);
not G5059 (W3662, W5051);
not G5060 (W3663, W5052);
not G5061 (W3664, W5053);
not G5062 (W3665, W5054);
not G5063 (W3666, W5055);
not G5064 (W3667, W5056);
not G5065 (W3668, W5057);
not G5066 (W3669, W5058);
not G5067 (W3670, W5059);
not G5068 (W3671, W5060);
not G5069 (W3672, W5061);
not G5070 (W3673, W5062);
not G5071 (W3674, W5063);
not G5072 (W3675, W5064);
not G5073 (W3676, W5065);
not G5074 (W3677, W5066);
not G5075 (W3678, W5067);
not G5076 (W3679, W5068);
not G5077 (W3680, W5069);
not G5078 (W3681, W5070);
not G5079 (W3682, W5071);
not G5080 (W3683, W5072);
not G5081 (W3684, W5073);
not G5082 (W3685, W5074);
not G5083 (W3686, W5075);
not G5084 (W3687, W5076);
not G5085 (W3688, W5077);
not G5086 (W3689, W5078);
not G5087 (W3690, W5079);
not G5088 (W3691, W5080);
not G5089 (W3692, W5081);
not G5090 (W3693, W5082);
not G5091 (W3694, W5083);
not G5092 (W3695, W5084);
not G5093 (W3696, W5085);
not G5094 (W3697, W5086);
not G5095 (W3698, W5087);
not G5096 (W3699, W5088);
not G5097 (W3700, W5089);
not G5098 (W3701, W5090);
not G5099 (W3702, W5091);
not G5100 (W3703, W5092);
not G5101 (W3704, W5093);
not G5102 (W3705, W5094);
not G5103 (W3706, W5095);
not G5104 (W3707, W5096);
not G5105 (W3708, W5097);
not G5106 (W3709, W5098);
not G5107 (W3710, W5099);
not G5108 (W3711, W5100);
not G5109 (W3712, W5101);
not G5110 (W3713, W5102);
not G5111 (W3714, W5103);
not G5112 (W3715, W5104);
not G5113 (W3716, W5105);
not G5114 (W3717, W5106);
not G5115 (W3718, W5107);
not G5116 (W3719, W5108);
not G5117 (W3720, W5109);
not G5118 (W3721, W5110);
not G5119 (W3722, W5111);
not G5120 (W3723, W5112);
not G5121 (W3724, W5113);
not G5122 (W3725, W5114);
not G5123 (W3726, W5115);
not G5124 (W3727, W5116);
not G5125 (W3728, W5117);
not G5126 (W3729, W5118);
not G5127 (W3730, W5119);
not G5128 (W3731, W5120);
not G5129 (W3732, W5121);
not G5130 (W3733, W5122);
not G5131 (W3734, W5123);
not G5132 (W3735, W5124);
not G5133 (W3736, W5125);
not G5134 (W3737, W5126);
not G5135 (W3738, W5127);
not G5136 (W3739, W5128);
not G5137 (W3740, W5129);
not G5138 (W3741, W5130);
not G5139 (W3742, W5131);
not G5140 (W3743, W5132);
not G5141 (W3744, W5133);
not G5142 (W3745, W5134);
not G5143 (W3746, W5135);
not G5144 (W3747, W5136);
not G5145 (W3748, W5137);
not G5146 (W3749, W5138);
not G5147 (W3750, W5139);
not G5148 (W3751, W5140);
not G5149 (W3752, W5141);
not G5150 (W3753, W5142);
not G5151 (W3754, W5143);
not G5152 (W3755, W5144);
not G5153 (W3756, W5145);
not G5154 (W3757, W5146);
not G5155 (W3758, W5147);
not G5156 (W3759, W5148);
not G5157 (W3760, W5149);
not G5158 (W3761, W5150);
not G5159 (W3762, W5151);
not G5160 (W3763, W5152);
not G5161 (W3764, W5153);
not G5162 (W3765, W5154);
not G5163 (W3766, W5155);
not G5164 (W3767, W5156);
not G5165 (W3768, W5157);
not G5166 (W3769, W5158);
not G5167 (W3770, W5159);
not G5168 (W3771, W5160);
not G5169 (W3772, W5161);
not G5170 (W3773, W5162);
not G5171 (W3774, W5163);
not G5172 (W3775, W5164);
not G5173 (W3776, W5165);
not G5174 (W3777, W5166);
not G5175 (W3778, W5167);
not G5176 (W3779, W5168);
not G5177 (W3780, W5169);
not G5178 (W3781, W5170);
not G5179 (W3782, W5171);
not G5180 (W3783, W5172);
not G5181 (W3784, W5173);
not G5182 (W3785, W5174);
not G5183 (W3786, W5175);
not G5184 (W3787, W5176);
not G5185 (W3788, W5177);
not G5186 (W3789, W5178);
not G5187 (W3790, W5179);
not G5188 (W3791, W5180);
not G5189 (W3792, W5181);
not G5190 (W3793, W5182);
not G5191 (W3794, W5183);
not G5192 (W3795, W5184);
not G5193 (W3796, W5185);
not G5194 (W3797, W5186);
not G5195 (W3798, W5187);
not G5196 (W3799, W5188);
not G5197 (W3800, W5189);
not G5198 (W3801, W5190);
not G5199 (W3802, W5191);
not G5200 (W3803, W5192);
not G5201 (W3804, W5193);
not G5202 (W3805, W5194);
not G5203 (W3806, W5195);
not G5204 (W3807, W5196);
not G5205 (W3808, W5197);
not G5206 (W3809, W5198);
not G5207 (W3810, W5199);
not G5208 (W3811, W5200);
not G5209 (W3812, W5201);
not G5210 (W3813, W5202);
not G5211 (W3814, W5203);
not G5212 (W3815, W5204);
not G5213 (W3816, W5205);
not G5214 (W3817, W5206);
not G5215 (W3818, W5207);
not G5216 (W3819, W5208);
not G5217 (W3820, W5209);
not G5218 (W3821, W5210);
not G5219 (W3822, W5211);
not G5220 (W3823, W5212);
not G5221 (W3824, W5213);
not G5222 (W3825, W5214);
not G5223 (W3826, W5215);
not G5224 (W3827, W5216);
not G5225 (W3828, W5217);
not G5226 (W3829, W5218);
not G5227 (W3830, W5219);
not G5228 (W3831, W5220);
not G5229 (W3832, W5221);
not G5230 (W3833, W5222);
not G5231 (W3834, W5223);
not G5232 (W3835, W5224);
not G5233 (W3836, W5225);
not G5234 (W3837, W5226);
not G5235 (W3838, W5227);
not G5236 (W3839, W5228);
not G5237 (W3840, W5229);
not G5238 (W3841, W5230);
not G5239 (W3842, W5231);
not G5240 (W3843, W5232);
not G5241 (W3844, W5233);
not G5242 (W3845, W5234);
not G5243 (W3846, W5235);
not G5244 (W3847, W5236);
not G5245 (W3848, W5237);
not G5246 (W3849, W5238);
not G5247 (W3850, W5239);
not G5248 (W3851, W5240);
not G5249 (W3852, W5241);
not G5250 (W3853, W5242);
not G5251 (W3854, W5243);
not G5252 (W3855, W5244);
not G5253 (W3856, W5245);
not G5254 (W3857, W5246);
not G5255 (W3858, W5247);
not G5256 (W3859, W5248);
not G5257 (W3860, W5249);
not G5258 (W3861, W5250);
not G5259 (W3862, W5251);
not G5260 (W3863, W5252);
not G5261 (W3864, W5253);
not G5262 (W3865, W5254);
not G5263 (W3866, W5255);
not G5264 (W3867, W5256);
not G5265 (W3868, W5257);
not G5266 (W3869, W5258);
not G5267 (W3870, W5259);
not G5268 (W3871, W5260);
not G5269 (W3872, W5261);
not G5270 (W3873, W5262);
not G5271 (W3874, W5263);
not G5272 (W3875, I222);
not G5273 (W3876, W5264);
not G5274 (W3877, W5265);
not G5275 (W3878, W5266);
not G5276 (W3879, W5267);
not G5277 (W3880, W5268);
not G5278 (W3881, W5269);
not G5279 (W3882, W5270);
not G5280 (W3883, W5271);
not G5281 (W3884, W5272);
not G5282 (W3885, W5273);
not G5283 (W3886, W5274);
not G5284 (W3887, W5275);
not G5285 (W3888, W5276);
not G5286 (W3889, W5277);
not G5287 (W3890, W5278);
not G5288 (W3891, W5279);
not G5289 (W3892, W5280);
not G5290 (W3893, W5281);
not G5291 (W3894, W5282);
not G5292 (W3895, W5283);
not G5293 (W3896, W5284);
not G5294 (W3897, W5285);
not G5295 (W3898, W5286);
not G5296 (W3899, W5287);
not G5297 (W3900, W5288);
not G5298 (W3901, W5289);
not G5299 (W3902, W5290);
not G5300 (W3903, W5291);
not G5301 (W3904, W5292);
not G5302 (W3905, W5293);
not G5303 (W3906, W5294);
not G5304 (W3907, W5295);
not G5305 (W3908, W5296);
not G5306 (W3909, W5297);
not G5307 (W3910, W5298);
not G5308 (W3911, W5299);
not G5309 (W3912, W5300);
not G5310 (W3913, W5301);
not G5311 (W3914, W5302);
not G5312 (W3915, W5303);
not G5313 (W3916, W5304);
not G5314 (W3917, W5305);
not G5315 (W3918, W5306);
not G5316 (W3919, W5307);
not G5317 (W3920, W5308);
not G5318 (W3921, W5309);
not G5319 (W3922, W5310);
not G5320 (W3923, W5311);
not G5321 (W3924, W5312);
not G5322 (W3925, W5313);
not G5323 (W3926, W5314);
not G5324 (W3927, W5315);
not G5325 (W3928, W5316);
not G5326 (W3929, W5317);
not G5327 (W3930, W5318);
not G5328 (W3931, W5319);
not G5329 (W3932, W5320);
not G5330 (W3933, W5321);
not G5331 (W3934, W5322);
not G5332 (W3935, W5323);
not G5333 (W3936, W5324);
not G5334 (W3937, W5325);
not G5335 (W3938, W5326);
not G5336 (W3939, W5327);
not G5337 (W3940, W5328);
not G5338 (W3941, W5329);
not G5339 (W3942, W5330);
not G5340 (W3943, W5331);
not G5341 (W3944, W5332);
not G5342 (W3945, W5333);
not G5343 (W3946, W5334);
not G5344 (W3947, W5335);
not G5345 (W3948, W5336);
not G5346 (W3949, W5337);
not G5347 (W3950, W5338);
not G5348 (W3951, W5339);
not G5349 (W3952, W5340);
not G5350 (W3953, W5341);
not G5351 (W3954, W5342);
not G5352 (W3955, W5343);
not G5353 (W3956, W5344);
not G5354 (W3957, W5345);
not G5355 (W3958, W5346);
not G5356 (W3959, W5347);
not G5357 (W3960, W5348);
not G5358 (W3961, W5349);
not G5359 (W3962, W5350);
not G5360 (W3963, W5351);
not G5361 (W3964, W5352);
not G5362 (W3965, W5353);
not G5363 (W3966, W5354);
not G5364 (W3967, W5355);
not G5365 (W3968, W5356);
not G5366 (W3969, W5357);
not G5367 (W3970, W5358);
not G5368 (W3971, W5359);
not G5369 (W3972, W5360);
not G5370 (W3973, W5361);
not G5371 (W3974, W5362);
not G5372 (W3975, W5363);
not G5373 (W3976, W5364);
not G5374 (W3977, W5365);
not G5375 (W3978, W5366);
not G5376 (W3979, W5367);
not G5377 (W3980, W5368);
not G5378 (W3981, W5369);
not G5379 (W3982, W5370);
not G5380 (W3983, W5371);
not G5381 (W3984, W5372);
not G5382 (W3985, W5373);
not G5383 (W3986, W5374);
not G5384 (W3987, W5375);
not G5385 (W3988, W5376);
not G5386 (W3989, W5377);
not G5387 (W3990, W5378);
not G5388 (W3991, W5379);
not G5389 (W3992, W5380);
not G5390 (W3993, W5381);
not G5391 (W3994, W5382);
not G5392 (W3995, W5383);
not G5393 (W3996, W5384);
not G5394 (W3997, W5385);
not G5395 (W3998, W5386);
not G5396 (W3999, W5387);
not G5397 (W4000, W5388);
not G5398 (W4001, W5389);
not G5399 (W4002, W5390);
not G5400 (W4003, W5391);
not G5401 (W4004, W5392);
not G5402 (W4005, W5393);
not G5403 (W4006, W5394);
not G5404 (W4007, W5395);
not G5405 (W4008, W5396);
not G5406 (W4009, W5397);
not G5407 (W4010, W5398);
not G5408 (W4011, W5399);
not G5409 (W4012, W5400);
not G5410 (W4013, W5401);
not G5411 (W4014, W5402);
not G5412 (W4015, W5403);
not G5413 (W4016, W5404);
not G5414 (W4017, W5405);
not G5415 (W4018, W5406);
not G5416 (W4019, W5407);
not G5417 (W4020, W5408);
not G5418 (W4021, W5409);
not G5419 (W4022, W5410);
not G5420 (W4023, W5411);
not G5421 (W4024, W5412);
not G5422 (W4025, W5413);
not G5423 (W4026, W5414);
not G5424 (W4027, W5415);
not G5425 (W4028, W5416);
not G5426 (W4029, W5417);
not G5427 (W4030, W5418);
not G5428 (W4031, W5419);
not G5429 (W4032, W5420);
not G5430 (W4033, W5421);
not G5431 (W4034, W5422);
not G5432 (W4035, W5423);
not G5433 (W4036, W5424);
not G5434 (W4037, W5425);
not G5435 (W4038, W5426);
not G5436 (W4039, W5427);
not G5437 (W4040, W5428);
not G5438 (W4041, W5429);
not G5439 (W4042, W5430);
not G5440 (W4043, W5431);
not G5441 (W4044, W5432);
not G5442 (W4045, W5433);
not G5443 (W4046, W5434);
not G5444 (W4047, W5435);
not G5445 (W4048, W5436);
not G5446 (W4049, W5437);
not G5447 (W4050, W5438);
not G5448 (W4051, W5439);
not G5449 (W4052, W5440);
not G5450 (W4053, W5441);
not G5451 (W4054, W5442);
not G5452 (W4055, W5443);
not G5453 (W4056, W5444);
not G5454 (W4057, W5445);
not G5455 (W4058, W5446);
not G5456 (W4059, W5447);
not G5457 (W4060, W5448);
not G5458 (W4061, W5449);
not G5459 (W4062, W5450);
not G5460 (W4063, W5451);
not G5461 (W4064, W5452);
not G5462 (W4065, W5453);
not G5463 (W4066, W5454);
not G5464 (W4067, W5455);
not G5465 (W4068, W5455);
not G5466 (W4069, W5455);
not G5467 (W4070, W5455);
not G5468 (W4071, W5455);
not G5469 (W4072, W5456);
not G5470 (W4073, W5456);
not G5471 (W4074, W5456);
not G5472 (W4075, W5456);
not G5473 (W4076, W5457);
not G5474 (W4077, W5458);
not G5475 (W4078, W5459);
not G5476 (W4079, W5460);
not G5477 (W4080, W5461);
not G5478 (W4081, W5461);
not G5479 (W4082, W5461);
not G5480 (W4083, W5462);
not G5481 (W4084, W5462);
not G5482 (W4085, W5463);
not G5483 (W4086, W5464);
not G5484 (W4087, W5464);
not G5485 (W4088, W5464);
not G5486 (W4089, W5465);
not G5487 (W4090, W5466);
not G5488 (W4091, W5467);
not G5489 (W4092, W5468);
not G5490 (W4093, W5469);
not G5491 (W4094, W5470);
not G5492 (W4095, W5471);
not G5493 (W4096, W5472);
not G5494 (W4097, W5473);
not G5495 (W4098, W5474);
not G5496 (W4099, W5475);
not G5497 (W4100, W5476);
not G5498 (W4101, W5477);
not G5499 (W4102, W5478);
not G5500 (W4103, W5479);
not G5501 (W4104, W5480);
not G5502 (W4105, W5481);
not G5503 (W4106, W5482);
not G5504 (W4107, W5483);
not G5505 (W4108, W5484);
not G5506 (W4109, W5485);
not G5507 (W4110, W5486);
not G5508 (W4111, W5487);
not G5509 (W4112, W5488);
not G5510 (W4113, W5489);
not G5511 (W4114, W5490);
not G5512 (W4115, W5491);
not G5513 (W4116, W5492);
not G5514 (W4117, W5493);
not G5515 (W4118, W5494);
not G5516 (W4119, W5495);
not G5517 (W4120, W5496);
not G5518 (W4121, W5497);
not G5519 (W4122, W5498);
not G5520 (W4123, W5499);
not G5521 (W4124, W5500);
not G5522 (W4125, W5501);
not G5523 (W4126, W5502);
not G5524 (W4127, W5503);
not G5525 (W4128, W5504);
not G5526 (W4129, W5505);
not G5527 (W4130, W5506);
not G5528 (W4131, W5507);
not G5529 (W4132, W5508);
not G5530 (W4133, W5509);
not G5531 (W4134, W5510);
not G5532 (W4135, W5511);
not G5533 (W4136, W5512);
not G5534 (W4137, W5513);
not G5535 (W4138, W5514);
not G5536 (W4139, W5515);
not G5537 (W4140, W5516);
not G5538 (W4141, W5517);
not G5539 (W4142, W5518);
not G5540 (W4143, W5519);
not G5541 (W4144, W5520);
not G5542 (W4145, W5521);
not G5543 (W4146, W5522);
not G5544 (W4147, W5523);
not G5545 (W4148, W5524);
not G5546 (W4149, W5525);
not G5547 (W4150, W5526);
not G5548 (W4151, W5527);
not G5549 (W4152, W5528);
not G5550 (W4153, W5529);
not G5551 (W4154, W5530);
not G5552 (W4155, W5531);
not G5553 (W4156, W5532);
not G5554 (W4157, W5533);
not G5555 (W4158, W5534);
not G5556 (W4159, W5535);
not G5557 (W4160, W5536);
not G5558 (W4161, W5537);
not G5559 (W4162, W5538);
not G5560 (W4163, W5539);
not G5561 (W4164, W5540);
not G5562 (W4165, W5541);
not G5563 (W4166, W5542);
not G5564 (W4167, W5543);
not G5565 (W4168, W5544);
not G5566 (W4169, W5545);
not G5567 (W4170, W5546);
not G5568 (W4171, W5547);
not G5569 (W4172, W5548);
not G5570 (W4173, W5549);
not G5571 (W4174, W5550);
not G5572 (W4175, W5551);
not G5573 (W4176, W5552);
not G5574 (W4177, W5553);
not G5575 (W4178, W5554);
not G5576 (W4179, W5555);
not G5577 (W4180, W5556);
not G5578 (W4181, W5557);
not G5579 (W4182, W5558);
not G5580 (W4183, W5559);
not G5581 (W4184, W5560);
not G5582 (W4185, W5561);
not G5583 (W4186, W5562);
not G5584 (W4187, W5563);
not G5585 (W4188, W5564);
not G5586 (W4189, W5565);
not G5587 (W4190, W5566);
not G5588 (W4191, W5567);
not G5589 (W4192, W5568);
not G5590 (W4193, W4192);
not G5591 (W4194, W5569);
not G5592 (W4195, W4194);
not G5593 (W4196, W4194);
not G5594 (W4197, W5570);
nand G5595 (W4198, W5571, W5572);
not G5596 (W4199, W5573);
nand G5597 (W4200, W5574, W5575);
nor G5598 (W4201, W5576, W5577);
nor G5599 (W4202, W5578, W5579);
nor G5600 (W4203, W5580, W5581);
nor G5601 (W4204, W5582, W5583);
nor G5602 (W4205, W5584, W5585);
nor G5603 (W4206, W5586, W5587);
nor G5604 (W4207, W5588, W5589);
nor G5605 (W4208, W5590, W5591);
nor G5606 (W4209, W5592, W5593);
nor G5607 (W4210, W5594, W5595);
nor G5608 (W4211, W5596, W5597);
nor G5609 (W4212, W5598, W5599);
nor G5610 (W4213, W5600, W5601);
nor G5611 (W4214, W5602, W5603);
nor G5612 (W4215, W5604, W5605);
nor G5613 (W4216, W5606, W5607);
nor G5614 (W4217, W5608, W5609);
nor G5615 (W4218, W5610, W5611);
nand G5616 (W4219, W5612, W5613);
nor G5617 (W4220, W5614, W5615);
nor G5618 (W4221, W5616, W5617);
nor G5619 (W4222, W5618, W5619);
nor G5620 (W4223, W5620, W5621);
nor G5621 (W4224, W5622, W5623);
nor G5622 (W4225, W5624, W5625);
nor G5623 (W4226, W5626, W5627);
nor G5624 (W4227, W5628, W5629);
nor G5625 (W4228, W5630, W5631);
nor G5626 (W4229, W5632, W5633);
nor G5627 (W4230, W5634, W5635);
nor G5628 (W4231, W5636, W5637);
nor G5629 (W4232, W5638, W5639);
nor G5630 (W4233, W5640, W5641);
nor G5631 (W4234, W5642, W5643);
nor G5632 (W4235, W5644, W5645);
nor G5633 (W4236, W5646, W5647);
nor G5634 (W4237, W5648, W5649);
nor G5635 (W4238, W5650, W5651);
nor G5636 (W4239, W5652, W5653);
nor G5637 (W4240, W5654, W5655);
nor G5638 (W4241, W5656, W5657);
nor G5639 (W4242, W5658, W5659);
nor G5640 (W4243, W5660, W5661);
nor G5641 (W4244, W5662, W5663);
nor G5642 (W4245, W5664, W5665);
nor G5643 (W4246, W5666, W5667);
nor G5644 (W4247, W5668, W5669);
nor G5645 (W4248, W5670, W5671);
nor G5646 (W4249, W5672, W5673);
nor G5647 (W4250, W5674, W5675);
nor G5648 (W4251, W5676, W5677);
nor G5649 (W4252, W5678, W5679);
nor G5650 (W4253, W5680, W5681);
nor G5651 (W4254, W5682, W5683);
nor G5652 (W4255, W5684, W5685);
nor G5653 (W4256, W5686, W5687);
nor G5654 (W4257, W5688, W5689);
nor G5655 (W4258, W5690, W5691);
nor G5656 (W4259, W5692, W5693);
nor G5657 (W4260, W5694, W5695);
nor G5658 (W4261, W5696, W5697);
nor G5659 (W4262, W5698, W5699);
nor G5660 (W4263, W5700, W5701);
nor G5661 (W4264, W5702, W5703);
nor G5662 (W4265, W5704, W5705);
nor G5663 (W4266, W5706, W5707);
nor G5664 (W4267, W5708, W5709);
nor G5665 (W4268, W5710, W5711);
nor G5666 (W4269, W5712, W5713);
nor G5667 (W4270, W5714, W5715);
nor G5668 (W4271, W5716, W5717);
nor G5669 (W4272, W5718, W5719);
nor G5670 (W4273, W5720, W5719);
nor G5671 (W4274, W5721, W5719);
nand G5672 (W4275, W5722, W5723);
nor G5673 (W4276, W5724, W5725);
nor G5674 (W4277, W5726, W5727);
nor G5675 (W4278, W5728, W5729);
nor G5676 (W4279, W5730, W5731);
nor G5677 (W4280, W5732, W5733);
nor G5678 (W4281, W5734, W5735);
nor G5679 (W4282, W5736, W5737);
nor G5680 (W4283, W5738, W5739);
nor G5681 (W4284, W5740, W5741);
nor G5682 (W4285, W5742, W5743);
nor G5683 (W4286, W5744, W5745);
nor G5684 (W4287, W5746, W5747);
nor G5685 (W4288, W5748, W5749);
nor G5686 (W4289, W5750, W5751);
nor G5687 (W4290, W5752, W5753);
nor G5688 (W4291, W5754, W5755);
nor G5689 (W4292, W5756, W5757);
nor G5690 (W4293, W5758, W5759);
nor G5691 (W4294, W5760, W5761);
nor G5692 (W4295, W5762, W5763);
nor G5693 (W4296, W5764, W5765);
nor G5694 (W4297, W5766, W5767);
nor G5695 (W4298, W5768, W5769);
nor G5696 (W4299, W5770, W5771);
nor G5697 (W4300, W5772, W5773);
nor G5698 (W4301, W5774, W5775);
nor G5699 (W4302, W5776, W5777);
nor G5700 (W4303, W5778, W5779);
nor G5701 (W4304, W5780, W5781);
nor G5702 (W4305, W5782, W5783);
nor G5703 (W4306, W5784, W5785);
nor G5704 (W4307, W5786, W5787);
nor G5705 (W4308, W5788, W5789);
nor G5706 (W4309, W5790, W5791);
nor G5707 (W4310, W5792, W5793);
nor G5708 (W4311, W5794, W5795);
nor G5709 (W4312, W5796, W5797);
nor G5710 (W4313, W5798, W5799);
nor G5711 (W4314, W5800, W5801);
nor G5712 (W4315, W5802, W5803);
nor G5713 (W4316, W5804, W5805);
nor G5714 (W4317, W5806, W5807);
nor G5715 (W4318, W5808, W5809);
nor G5716 (W4319, W5810, W5811);
nor G5717 (W4320, W5812, W5813);
nor G5718 (W4321, W5814, W5815);
nor G5719 (W4322, W5816, W5817);
nor G5720 (W4323, W5818, W5819);
nor G5721 (W4324, W5820, W5821);
nor G5722 (W4325, W5822, W5823);
nor G5723 (W4326, W5824, W5825);
nor G5724 (W4327, W5826, W5827);
nor G5725 (W4328, W5828, W5829);
nor G5726 (W4329, W5830, W5831);
nor G5727 (W4330, W5832, W5833);
nor G5728 (W4331, W5834, W5835);
nor G5729 (W4332, W5836, W5837);
nor G5730 (W4333, W5838, W5839);
nor G5731 (W4334, W5840, W5841);
nor G5732 (W4335, W5842, W5837);
nor G5733 (W4336, W5843, W5837);
nor G5734 (W4337, W5844, W5837);
nor G5735 (W4338, W5845, W5837);
nor G5736 (W4339, W5846, W5847);
not G5737 (W4340, W5848);
not G5738 (W4341, W5849);
not G5739 (W4342, W5850);
not G5740 (W4343, W5851);
not G5741 (W4344, W5852);
not G5742 (W4345, W5853);
not G5743 (W4346, W5854);
not G5744 (W4347, W5855);
not G5745 (W4348, W5856);
not G5746 (W4349, W5857);
not G5747 (W4350, W5858);
not G5748 (W4351, W5859);
not G5749 (W4352, W5860);
nand G5750 (W4353, W5861, W5862);
nor G5751 (W4354, W5863, W5847);
not G5752 (W4355, W5864);
not G5753 (W4356, W5865);
not G5754 (W4357, W5866);
not G5755 (W4358, W5867);
not G5756 (W4359, W5868);
not G5757 (W4360, W5869);
not G5758 (W4361, W5870);
not G5759 (W4362, W5871);
not G5760 (W4363, W5872);
nor G5761 (W4364, W5873, W5874);
nor G5762 (W4365, W5875, W5876);
nor G5763 (W4366, W5877, W5878);
nor G5764 (W4367, W5879, W5880);
nor G5765 (W4368, W5881, W5882);
nor G5766 (W4369, W5883, W5884);
nor G5767 (W4370, W5885, W5886);
nor G5768 (W4371, W5887, W5888);
nor G5769 (W4372, W5889, W5890);
nor G5770 (W4373, W5891, W5892);
nor G5771 (W4374, W5893, W5894);
nor G5772 (W4375, W5895, W5896);
nor G5773 (W4376, W5897, W5898);
nor G5774 (W4377, W5899, W5900);
nor G5775 (W4378, W5901, W5902);
nor G5776 (W4379, W5903, W5904);
nor G5777 (W4380, W5905, W5906);
nor G5778 (W4381, W5907, W5908);
nor G5779 (W4382, W5909, W5910);
nor G5780 (W4383, W5911, W5912);
nor G5781 (W4384, W5913, W5914);
nor G5782 (W4385, W5915, W5916);
nor G5783 (W4386, W5917, W5918);
nor G5784 (W4387, W5919, W5920);
nor G5785 (W4388, W5921, W5922);
nor G5786 (W4389, W5923, W5924);
nor G5787 (W4390, W5925, W5926);
nor G5788 (W4391, W5927, W5928);
nor G5789 (W4392, W5929, W5930);
nor G5790 (W4393, W5931, W5932);
nor G5791 (W4394, W5933, W5934);
nor G5792 (W4395, W5935, W5936);
nor G5793 (W4396, W5937, W5938);
nor G5794 (W4397, W5939, W5940);
nor G5795 (W4398, W5941, W5942);
nor G5796 (W4399, W5943, W5944);
nor G5797 (W4400, W5945, W5946);
nor G5798 (W4401, W5947, W5948);
nor G5799 (W4402, W5949, W5950);
nor G5800 (W4403, W5951, W5952);
nor G5801 (W4404, W5953, W5954);
nor G5802 (W4405, W5955, W5956);
nor G5803 (W4406, W5957, W5958);
nor G5804 (W4407, W5959, W5958);
nor G5805 (W4408, W5960, W5958);
nor G5806 (W4409, W5961, W5958);
nor G5807 (W4410, W5962, W5958);
nor G5808 (W4411, W5963, W5958);
nor G5809 (W4412, W5964, W5958);
nor G5810 (W4413, W5965, W5958);
nor G5811 (W4414, W5966, W5958);
nor G5812 (W4415, W5967, W5958);
nor G5813 (W4416, W5968, W5969);
nor G5814 (W4417, W5970, W5971);
nor G5815 (W4418, W5972, W5973);
nor G5816 (W4419, W5974, W5975);
nor G5817 (W4420, W5976, W5977);
nor G5818 (W4421, W5978, W5979);
nor G5819 (W4422, W5980, W5981);
nor G5820 (W4423, W5982, W5983);
nor G5821 (W4424, W5984, W5985);
not G5822 (W4425, W5986);
not G5823 (W4426, W5987);
not G5824 (W4427, W5988);
not G5825 (W4428, W5989);
nor G5826 (W4429, W5990, W5991);
nor G5827 (W4430, W5992, W5993);
nor G5828 (W4431, W5994, W5995);
nor G5829 (W4432, W5996, W5997);
nor G5830 (W4433, W5998, W5999);
nor G5831 (W4434, W6000, W6001);
nor G5832 (W4435, W6002, W6003);
nor G5833 (W4436, W6004, W6005);
nor G5834 (W4437, W6006, W6007);
nor G5835 (W4438, W6008, W6009);
not G5836 (W4439, W6010);
nor G5837 (W4440, W6011, W6012);
not G5838 (W4441, W6013);
nor G5839 (W4442, W6014, W6015);
not G5840 (W4443, W6016);
nor G5841 (W4444, W6017, W6018);
not G5842 (W4445, W6019);
nor G5843 (W4446, W6020, W6021);
nor G5844 (W4447, W6022, W6023);
nor G5845 (W4448, W6024, W6025);
not G5846 (W4449, W6026);
nor G5847 (W4450, W6027, W6028);
nor G5848 (W4451, W6029, W6030);
nor G5849 (W4452, W6031, W6032);
not G5850 (W4453, W6033);
nor G5851 (W4454, W6034, W6035);
not G5852 (W4455, W6036);
nor G5853 (W4456, W6037, W6038);
nor G5854 (W4457, W6039, W6040);
not G5855 (W4458, W6041);
not G5856 (W4459, W6042);
nor G5857 (W4460, W6043, W6044);
nor G5858 (W4461, W6045, W6046);
nor G5859 (W4462, W6047, W6048);
nor G5860 (W4463, W6049, W6050, W6051);
nor G5861 (W4464, W6052, W6053, W6054);
nor G5862 (W4465, W6055, W6056);
nor G5863 (W4466, W6057, W6058);
nor G5864 (W4467, W6059, W6060);
nor G5865 (W4468, W6061, W6062);
nor G5866 (W4469, W6063, W6064);
nor G5867 (W4470, W6065, W6066);
nor G5868 (W4471, W6067, W6068);
nor G5869 (W4472, W6069, W6070);
not G5870 (W4473, W6071);
not G5871 (W4474, W6072);
not G5872 (W4475, W6073);
not G5873 (W4476, W6074);
not G5874 (W4477, W6075);
not G5875 (W4478, W6076);
not G5876 (W4479, W6077);
not G5877 (W4480, W6078);
not G5878 (W4481, W6079);
not G5879 (W4482, W6080);
nor G5880 (W4483, W6081, W6082);
nor G5881 (W4484, W6083, W6084);
nor G5882 (W4485, W6085, W6086);
nor G5883 (W4486, W6087, W6088);
nor G5884 (W4487, W6089, W6090);
nor G5885 (W4488, W6091, W6092);
nor G5886 (W4489, W6093, W6094);
nor G5887 (W4490, W6095, W6096);
nor G5888 (W4491, W6097, W6098);
nor G5889 (W4492, W6099, W6100);
nor G5890 (W4493, W6101, W6102);
nor G5891 (W4494, W6103, W6104);
nor G5892 (W4495, W6105, W6106);
nor G5893 (W4496, W6107, W6108);
nor G5894 (W4497, W6109, W6110);
nor G5895 (W4498, W6111, W6112);
nor G5896 (W4499, W6113, W6114);
nor G5897 (W4500, W6115, W6116);
nor G5898 (W4501, W6117, W6118);
nor G5899 (W4502, W6119, W6120);
nor G5900 (W4503, W6121, W6122);
nor G5901 (W4504, W6123, W6124);
nor G5902 (W4505, W6125, W6126);
nor G5903 (W4506, W6127, W6128);
nor G5904 (W4507, W6129, W6130);
nor G5905 (W4508, W6131, W6132);
nor G5906 (W4509, W6133, W6134);
nor G5907 (W4510, W6135, W6136);
nor G5908 (W4511, W6137, W6138);
nor G5909 (W4512, W6139, W6140);
nor G5910 (W4513, W6141, W6142);
nor G5911 (W4514, W6143, W6144);
nor G5912 (W4515, W6145, W6146);
nor G5913 (W4516, W6147, W6148);
nor G5914 (W4517, W6149, W6150);
nor G5915 (W4518, W6151, W6152);
nor G5916 (W4519, W6153, W6154);
nor G5917 (W4520, W6155, W6156);
nor G5918 (W4521, W6157, W6158);
nor G5919 (W4522, W6159, W6160);
nor G5920 (W4523, W6161, W6162);
nor G5921 (W4524, W6163, W6164);
nor G5922 (W4525, W6165, W6166);
nor G5923 (W4526, W6167, W6168);
nor G5924 (W4527, W6169, W6170);
nand G5925 (W4528, W4529, W6171);
not G5926 (W4529, W6172);
nor G5927 (W4530, W6173, W6174);
nor G5928 (W4531, W6175, W6176);
nor G5929 (W4532, W6177, W6178);
nor G5930 (W4533, W6179, W6180);
nor G5931 (W4534, W6181, W6182);
nor G5932 (W4535, W6183, W6184);
nor G5933 (W4536, W6185, W6186);
nor G5934 (W4537, W6187, W6188);
nor G5935 (W4538, W6189, W6190);
nor G5936 (W4539, W6191, W6192);
nor G5937 (W4540, W6193, W6194);
nor G5938 (W4541, W6195, W6196);
nor G5939 (W4542, W6197, W6198);
nor G5940 (W4543, W6199, W6200);
nor G5941 (W4544, W6201, W6202);
nor G5942 (W4545, W6203, W6204);
nor G5943 (W4546, W6205, W6206);
nor G5944 (W4547, W6207, W6208);
nor G5945 (W4548, W6209, W6210);
nor G5946 (W4549, W6211, W6212);
nor G5947 (W4550, W6213, W6214);
nor G5948 (W4551, W6215, W6216);
nor G5949 (W4552, W6217, W6218);
nor G5950 (W4553, W6219, W6220);
nor G5951 (W4554, W6221, W6222);
nor G5952 (W4555, W6223, W6224);
nor G5953 (W4556, W6225, W6226);
nor G5954 (W4557, W6227, W6228);
nor G5955 (W4558, W6229, W6230);
nor G5956 (W4559, W6231, W6232);
not G5957 (W4560, W6233);
not G5958 (W4561, W6234);
not G5959 (W4562, W6235);
not G5960 (W4563, W6236);
not G5961 (W4564, W6237);
not G5962 (W4565, W6238);
not G5963 (W4566, W6239);
not G5964 (W4567, W6240);
not G5965 (W4568, W6241);
not G5966 (W4569, W6242);
not G5967 (W4570, W6243);
not G5968 (W4571, W6244);
not G5969 (W4572, W6245);
not G5970 (W4573, W6246);
not G5971 (W4574, W6247);
not G5972 (W4575, W6248);
not G5973 (W4576, W6249);
nor G5974 (W4577, W6250, W6251);
nor G5975 (W4578, W6252, W6253);
nor G5976 (W4579, W6254, W6255);
nor G5977 (W4580, W6256, W6257);
nor G5978 (W4581, W6258, W6259);
nor G5979 (W4582, W6260, W6261);
nor G5980 (W4583, W6262, W6263);
nor G5981 (W4584, W6264, W6265);
nor G5982 (W4585, W6266, W6267);
nor G5983 (W4586, W6268, W6269);
nor G5984 (W4587, W6270, W6271);
nor G5985 (W4588, W6272, W6273);
nor G5986 (W4589, W6274, W6275);
nor G5987 (W4590, W6276, W6277);
nor G5988 (W4591, W6278, W6279);
nor G5989 (W4592, W6280, W6281);
nor G5990 (W4593, W6282, W6283);
nor G5991 (W4594, W6284, W6285);
nor G5992 (W4595, W6286, W6287);
nor G5993 (W4596, W6288, W6289);
nor G5994 (W4597, W6290, W6291);
nor G5995 (W4598, W6292, W6293);
nor G5996 (W4599, W6294, W6295);
nor G5997 (W4600, W6296, W6297);
nor G5998 (W4601, W6298, W6299);
nor G5999 (W4602, W6300, W6301);
nor G6000 (W4603, W6302, W6303);
nor G6001 (W4604, W6304, W6305);
nor G6002 (W4605, W6306, W6307);
nor G6003 (W4606, W6308, W6309);
nor G6004 (W4607, W6310, W6311);
nor G6005 (W4608, W6312, W6311);
nor G6006 (W4609, W6313, W6311);
nor G6007 (W4610, W6314, W6311);
nor G6008 (W4611, W6315, W6311);
nor G6009 (W4612, W6316, W6311);
nor G6010 (W4613, W6317, W6311);
nor G6011 (W4614, W6318, W6311);
nor G6012 (W4615, W6319, W6311);
nor G6013 (W4616, W6320, W6311);
not G6014 (W4617, W6321);
nor G6015 (W4618, W6322, W6323);
nor G6016 (W4619, W6324, W6325);
nor G6017 (W4620, W6326, W6327);
nor G6018 (W4621, W6328, W6329);
nor G6019 (W4622, W6330, W6331);
nor G6020 (W4623, W6332, W6333);
nor G6021 (W4624, W6334, W6335);
nor G6022 (W4625, W6336, W6337);
nor G6023 (W4626, W6338, W6339);
nor G6024 (W4627, W6340, W6341);
nor G6025 (W4628, W6342, W6343);
nor G6026 (W4629, W6344, W6345);
not G6027 (W4630, W6346);
not G6028 (W4631, W6347);
not G6029 (W4632, W6348);
not G6030 (W4633, W6349);
not G6031 (W4634, W6350);
not G6032 (W4635, W6351);
not G6033 (W4636, W6352);
not G6034 (W4637, W6353);
not G6035 (W4638, W6354);
nor G6036 (W4639, W6355, W6356);
nor G6037 (W4640, W6357, W6358);
nor G6038 (W4641, W6359, W6360);
nor G6039 (W4642, W6361, W6362);
nor G6040 (W4643, W6363, W6364);
nor G6041 (W4644, W6365, W6366);
nor G6042 (W4645, W6367, W6368);
nor G6043 (W4646, W6369, W6370);
nor G6044 (W4647, W6371, W6372);
nor G6045 (W4648, W6373, W6374);
nor G6046 (W4649, W6375, W6376);
nor G6047 (W4650, W6377, W6378);
nor G6048 (W4651, W6379, W6380);
nor G6049 (W4652, W6381, W6382);
nor G6050 (W4653, W6383, W6384);
nor G6051 (W4654, W6385, W6386);
nor G6052 (W4655, W6387, W6388);
nor G6053 (W4656, W6389, W6390);
nor G6054 (W4657, W6391, W6392);
nor G6055 (W4658, W6393, W6394);
nor G6056 (W4659, W6395, W6396);
nor G6057 (W4660, W6397, W6398);
nor G6058 (W4661, W6399, W6400);
nor G6059 (W4662, W6401, W6402);
nor G6060 (W4663, W6403, W6404);
nor G6061 (W4664, W6405, W6406);
nor G6062 (W4665, W6407, W6408);
nor G6063 (W4666, W6409, W6410);
nor G6064 (W4667, W6411, W6412);
nor G6065 (W4668, W6413, W6414);
nor G6066 (W4669, W6415, W6416);
nor G6067 (W4670, W6417, W6418);
nor G6068 (W4671, W6419, W6420);
nor G6069 (W4672, W6421, W6422);
nor G6070 (W4673, W6423, W6424);
nor G6071 (W4674, W6425, W6426);
nor G6072 (W4675, W6427, W6428);
nor G6073 (W4676, W6429, W6430);
nor G6074 (W4677, W6431, W6432);
nor G6075 (W4678, W6433, W6434);
nor G6076 (W4679, W6435, W6436);
nor G6077 (W4680, W6437, W6438);
nor G6078 (W4681, W6439, W6440);
nor G6079 (W4682, W6441, W6440);
nor G6080 (W4683, W6442, W6440);
nor G6081 (W4684, W6443, W6440);
nor G6082 (W4685, W6444, W6440);
nor G6083 (W4686, W6445, W6440);
nor G6084 (W4687, W6446, W6440);
nor G6085 (W4688, W6447, W6440);
nor G6086 (W4689, W6448, W6440);
nor G6087 (W4690, W6449, W6440);
nor G6088 (W4691, W6450, W6451);
nor G6089 (W4692, W6452, W6453);
nor G6090 (W4693, W6454, W6455);
nor G6091 (W4694, W6456, W6457);
nor G6092 (W4695, W6458, W6459);
nor G6093 (W4696, W6460, W6461);
nor G6094 (W4697, W6462, W6463);
nor G6095 (W4698, W6464, W6465);
nor G6096 (W4699, W6466, W6467);
not G6097 (W4700, W6468);
not G6098 (W4701, W6469);
not G6099 (W4702, W6470);
not G6100 (W4703, W6471);
nor G6101 (W4704, W6472, W6473);
nor G6102 (W4705, W6474, W6475);
nor G6103 (W4706, W6476, W6477);
nor G6104 (W4707, W6478, W6479);
nor G6105 (W4708, W6480, W6481);
nor G6106 (W4709, W6482, W6483);
nor G6107 (W4710, W6484, W6485);
nor G6108 (W4711, W6486, W6487);
nor G6109 (W4712, W6488, W6489);
nor G6110 (W4713, W6490, W6491);
not G6111 (W4714, W6492);
nor G6112 (W4715, W6493, W6494);
not G6113 (W4716, W6495);
nor G6114 (W4717, W6496, W6497);
not G6115 (W4718, W6498);
nor G6116 (W4719, W6499, W6500);
not G6117 (W4720, W6501);
nor G6118 (W4721, W6502, W6503);
nor G6119 (W4722, W6504, W6505);
nor G6120 (W4723, W6506, W6507);
not G6121 (W4724, W6508);
nor G6122 (W4725, W6509, W6510);
nor G6123 (W4726, W6511, W6512);
nor G6124 (W4727, W6513, W6514);
not G6125 (W4728, W6515);
nor G6126 (W4729, W6516, W6517);
not G6127 (W4730, W6518);
nor G6128 (W4731, W6519, W6520);
nor G6129 (W4732, W6521, W6522);
not G6130 (W4733, W6523);
not G6131 (W4734, W6524);
nor G6132 (W4735, W6525, W6526);
nor G6133 (W4736, W6527, W6528);
nor G6134 (W4737, W6529, W6530);
nor G6135 (W4738, W6531, W6532, W6533);
nor G6136 (W4739, W6534, W6535, W6536);
nor G6137 (W4740, W6537, W6538);
nor G6138 (W4741, W6539, W6540);
nor G6139 (W4742, W6541, W6542);
nor G6140 (W4743, W6543, W6544);
nor G6141 (W4744, W6545, W6546);
nor G6142 (W4745, W6547, W6548);
nor G6143 (W4746, W6549, W6550);
nor G6144 (W4747, W6551, W6552);
not G6145 (W4748, W6553);
not G6146 (W4749, W6554);
not G6147 (W4750, W6555);
not G6148 (W4751, W6556);
not G6149 (W4752, W6557);
not G6150 (W4753, W6558);
not G6151 (W4754, W6559);
not G6152 (W4755, W6560);
not G6153 (W4756, W6561);
not G6154 (W4757, W6562);
nor G6155 (W4758, W6563, W6564);
nor G6156 (W4759, W6565, W6566);
nor G6157 (W4760, W6567, W6568);
nor G6158 (W4761, W6569, W6570);
nor G6159 (W4762, W6571, W6572);
nor G6160 (W4763, W6573, W6574);
nor G6161 (W4764, W6575, W6576);
nor G6162 (W4765, W6577, W6578);
nor G6163 (W4766, W6579, W6580);
nor G6164 (W4767, W6581, W6582);
nor G6165 (W4768, W6583, W6584);
nor G6166 (W4769, W6585, W6586);
nor G6167 (W4770, W6587, W6588);
nor G6168 (W4771, W6589, W6590);
nor G6169 (W4772, W6591, W6592);
nor G6170 (W4773, W6593, W6594);
nor G6171 (W4774, W6595, W6596);
nor G6172 (W4775, W6597, W6598);
nor G6173 (W4776, W6599, W6600);
nor G6174 (W4777, W6601, W6602);
nor G6175 (W4778, W6603, W6604);
nor G6176 (W4779, W6605, W6606);
nor G6177 (W4780, W6607, W6608);
nor G6178 (W4781, W6609, W6610);
nor G6179 (W4782, W6611, W6612);
nor G6180 (W4783, W6613, W6614);
nor G6181 (W4784, W6615, W6616);
nor G6182 (W4785, W6617, W6618);
nor G6183 (W4786, W6619, W6620);
nor G6184 (W4787, W6621, W6622);
nor G6185 (W4788, W6623, W6624);
nor G6186 (W4789, W6625, W6626);
nor G6187 (W4790, W6627, W6628);
nor G6188 (W4791, W6629, W6630);
nor G6189 (W4792, W6631, W6632);
nor G6190 (W4793, W6633, W6634);
nor G6191 (W4794, W6635, W6636);
nor G6192 (W4795, W6637, W6638);
nor G6193 (W4796, W6639, W6640);
nor G6194 (W4797, W6641, W6642);
nor G6195 (W4798, W6643, W6644);
nor G6196 (W4799, W6645, W6646);
nor G6197 (W4800, W6647, W6648);
nor G6198 (W4801, W6649, W6650);
nor G6199 (W4802, W6651, W6652);
nand G6200 (W4803, W4804, W6653);
not G6201 (W4804, W6654);
nor G6202 (W4805, W6655, W6656);
nor G6203 (W4806, W6657, W6658);
nor G6204 (W4807, W6659, W6660);
nor G6205 (W4808, W6661, W6662);
nor G6206 (W4809, W6663, W6664);
nor G6207 (W4810, W6665, W6666);
nor G6208 (W4811, W6667, W6668);
nor G6209 (W4812, W6669, W6670);
nor G6210 (W4813, W6671, W6672);
nor G6211 (W4814, W6673, W6674);
nor G6212 (W4815, W6675, W6676);
nor G6213 (W4816, W6677, W6678);
nor G6214 (W4817, W6679, W6680);
nor G6215 (W4818, W6681, W6682);
nor G6216 (W4819, W6683, W6684);
nor G6217 (W4820, W6685, W6686);
nor G6218 (W4821, W6687, W6688);
nor G6219 (W4822, W6689, W6690);
nor G6220 (W4823, W6691, W6692);
nor G6221 (W4824, W6693, W6694);
nor G6222 (W4825, W6695, W6696);
nor G6223 (W4826, W6697, W6698);
nor G6224 (W4827, W6699, W6700);
nor G6225 (W4828, W6701, W6702);
nor G6226 (W4829, W6703, W6704);
nor G6227 (W4830, W6705, W6706);
nor G6228 (W4831, W6707, W6708);
nor G6229 (W4832, W6709, W6710);
nor G6230 (W4833, W6711, W6712);
nor G6231 (W4834, W6713, W6714);
not G6232 (W4835, W6715);
not G6233 (W4836, W6716);
not G6234 (W4837, W6717);
not G6235 (W4838, W6718);
not G6236 (W4839, W6719);
not G6237 (W4840, W6720);
not G6238 (W4841, W6721);
not G6239 (W4842, W6722);
not G6240 (W4843, W6723);
not G6241 (W4844, W6724);
not G6242 (W4845, W6725);
not G6243 (W4846, W6726);
not G6244 (W4847, W6727);
not G6245 (W4848, W6728);
not G6246 (W4849, W6729);
not G6247 (W4850, W6730);
not G6248 (W4851, W6731);
nor G6249 (W4852, W6732, W6733);
nor G6250 (W4853, W6734, W6735);
nor G6251 (W4854, W6736, W6737);
nor G6252 (W4855, W6738, W6739);
nor G6253 (W4856, W6740, W6741);
nor G6254 (W4857, W6742, W6743);
nor G6255 (W4858, W6744, W6745);
nor G6256 (W4859, W6746, W6747);
nor G6257 (W4860, W6748, W6749);
nor G6258 (W4861, W6750, W6751);
nor G6259 (W4862, W6752, W6753);
nor G6260 (W4863, W6754, W6755);
nor G6261 (W4864, W6756, W6757);
nor G6262 (W4865, W6758, W6759);
nor G6263 (W4866, W6760, W6761);
nor G6264 (W4867, W6762, W6763);
nor G6265 (W4868, W6764, W6765);
nor G6266 (W4869, W6766, W6767);
nor G6267 (W4870, W6768, W6769);
nor G6268 (W4871, W6770, W6771);
nor G6269 (W4872, W6772, W6773);
nor G6270 (W4873, W6774, W6775);
nor G6271 (W4874, W6776, W6777);
nor G6272 (W4875, W6778, W6779);
nor G6273 (W4876, W6780, W6781);
nor G6274 (W4877, W6782, W6783);
nor G6275 (W4878, W6784, W6785);
nor G6276 (W4879, W6786, W6787);
nor G6277 (W4880, W6788, W6789);
nor G6278 (W4881, W6790, W6791);
nor G6279 (W4882, W6792, W6793);
nor G6280 (W4883, W6794, W6793);
nor G6281 (W4884, W6795, W6793);
nor G6282 (W4885, W6796, W6793);
nor G6283 (W4886, W6797, W6793);
nor G6284 (W4887, W6798, W6793);
nor G6285 (W4888, W6799, W6793);
nor G6286 (W4889, W6800, W6793);
nor G6287 (W4890, W6801, W6793);
nor G6288 (W4891, W6802, W6793);
not G6289 (W4892, W6803);
nor G6290 (W4893, W6804, W6805);
nor G6291 (W4894, W6806, W6807);
nor G6292 (W4895, W6808, W6809);
nor G6293 (W4896, W6810, W6811);
nor G6294 (W4897, W6812, W6813);
nor G6295 (W4898, W6814, W6815);
nor G6296 (W4899, W6816, W6817);
nor G6297 (W4900, W6818, W6819);
nor G6298 (W4901, W6820, W6821);
nor G6299 (W4902, W6822, W6823);
nor G6300 (W4903, W6824, W6825);
nor G6301 (W4904, W6826, W6827);
not G6302 (W4905, W6828);
not G6303 (W4906, W6829);
not G6304 (W4907, W6830);
not G6305 (W4908, W6831);
not G6306 (W4909, W6832);
not G6307 (W4910, W6833);
not G6308 (W4911, W6834);
not G6309 (W4912, W6835);
not G6310 (W4913, W6836);
nor G6311 (W4914, W6837, W6838);
nor G6312 (W4915, W6839, W6840);
nor G6313 (W4916, W6841, W6842);
nor G6314 (W4917, W6843, W6844);
nor G6315 (W4918, W6845, W6846);
nor G6316 (W4919, W6847, W6848);
nor G6317 (W4920, W6849, W6850);
nor G6318 (W4921, W6851, W6852);
nor G6319 (W4922, W6853, W6854);
nor G6320 (W4923, W6855, W6856);
nor G6321 (W4924, W6857, W6858);
nor G6322 (W4925, W6859, W6860);
nor G6323 (W4926, W6861, W6862);
nor G6324 (W4927, W6863, W6864);
nor G6325 (W4928, W6865, W6866);
nor G6326 (W4929, W6867, W6868);
nor G6327 (W4930, W6869, W6870);
nor G6328 (W4931, W6871, W6872);
nor G6329 (W4932, W6873, W6874);
nor G6330 (W4933, W6875, W6876);
nor G6331 (W4934, W6877, W6878);
nor G6332 (W4935, W6879, W6880);
nor G6333 (W4936, W6881, W6882);
nor G6334 (W4937, W6883, W6884);
nor G6335 (W4938, W6885, W6886);
nor G6336 (W4939, W6887, W6888);
nor G6337 (W4940, W6889, W6890);
nor G6338 (W4941, W6891, W6892);
nor G6339 (W4942, W6893, W6894);
nor G6340 (W4943, W6895, W6896);
nor G6341 (W4944, W6897, W6898);
nor G6342 (W4945, W6899, W6900);
nor G6343 (W4946, W6901, W6902);
nor G6344 (W4947, W6903, W6904);
nor G6345 (W4948, W6905, W6906);
nor G6346 (W4949, W6907, W6908);
nor G6347 (W4950, W6909, W6910);
nor G6348 (W4951, W6911, W6912);
nor G6349 (W4952, W6913, W6914);
nor G6350 (W4953, W6915, W6916);
nor G6351 (W4954, W6917, W6918);
nor G6352 (W4955, W6919, W6920);
nor G6353 (W4956, W6921, W6922);
nor G6354 (W4957, W6923, W6922);
nor G6355 (W4958, W6924, W6922);
nor G6356 (W4959, W6925, W6922);
nor G6357 (W4960, W6926, W6922);
nor G6358 (W4961, W6927, W6922);
nor G6359 (W4962, W6928, W6922);
nor G6360 (W4963, W6929, W6922);
nor G6361 (W4964, W6930, W6922);
nor G6362 (W4965, W6931, W6922);
nor G6363 (W4966, W6932, W6933);
nor G6364 (W4967, W6934, W6935);
nor G6365 (W4968, W6936, W6937);
nor G6366 (W4969, W6938, W6939);
nor G6367 (W4970, W6940, W6941);
nor G6368 (W4971, W6942, W6943);
nor G6369 (W4972, W6944, W6945);
nor G6370 (W4973, W6946, W6947);
nor G6371 (W4974, W6948, W6949);
not G6372 (W4975, W6950);
not G6373 (W4976, W6951);
not G6374 (W4977, W6952);
not G6375 (W4978, W6953);
nor G6376 (W4979, W6954, W6955);
nor G6377 (W4980, W6956, W6957);
nor G6378 (W4981, W6958, W6959);
nor G6379 (W4982, W6960, W6961);
nor G6380 (W4983, W6962, W6963);
nor G6381 (W4984, W6964, W6965);
nor G6382 (W4985, W6966, W6967);
nor G6383 (W4986, W6968, W6969);
nor G6384 (W4987, W6970, W6971);
nor G6385 (W4988, W6972, W6973);
not G6386 (W4989, W6974);
nor G6387 (W4990, W6975, W6976);
not G6388 (W4991, W6977);
nor G6389 (W4992, W6978, W6979);
not G6390 (W4993, W6980);
nor G6391 (W4994, W6981, W6982);
not G6392 (W4995, W6983);
nor G6393 (W4996, W6984, W6985);
nor G6394 (W4997, W6986, W6987);
nor G6395 (W4998, W6988, W6989);
not G6396 (W4999, W6990);
nor G6397 (W5000, W6991, W6992);
nor G6398 (W5001, W6993, W6994);
nor G6399 (W5002, W6995, W6996);
not G6400 (W5003, W6997);
nor G6401 (W5004, W6998, W6999);
not G6402 (W5005, W7000);
nor G6403 (W5006, W7001, W7002);
nor G6404 (W5007, W7003, W7004);
not G6405 (W5008, W7005);
not G6406 (W5009, W7006);
nor G6407 (W5010, W7007, W7008);
nor G6408 (W5011, W7009, W7010);
nor G6409 (W5012, W7011, W7012);
nor G6410 (W5013, W7013, W7014, W7015);
nor G6411 (W5014, W7016, W7017, W7018);
nor G6412 (W5015, W7019, W7020);
nor G6413 (W5016, W7021, W7022);
nor G6414 (W5017, W7023, W7024);
nor G6415 (W5018, W7025, W7026);
nor G6416 (W5019, W7027, W7028);
nor G6417 (W5020, W7029, W7030);
nor G6418 (W5021, W7031, W7032);
nor G6419 (W5022, W7033, W7034);
not G6420 (W5023, W7035);
not G6421 (W5024, W7036);
not G6422 (W5025, W7037);
not G6423 (W5026, W7038);
not G6424 (W5027, W7039);
not G6425 (W5028, W7040);
not G6426 (W5029, W7041);
not G6427 (W5030, W7042);
not G6428 (W5031, W7043);
not G6429 (W5032, W7044);
nor G6430 (W5033, W7045, W7046);
nor G6431 (W5034, W7047, W7048);
nor G6432 (W5035, W7049, W7050);
nor G6433 (W5036, W7051, W7052);
nor G6434 (W5037, W7053, W7054);
nor G6435 (W5038, W7055, W7056);
nor G6436 (W5039, W7057, W7058);
nor G6437 (W5040, W7059, W7060);
nor G6438 (W5041, W7061, W7062);
nor G6439 (W5042, W7063, W7064);
nor G6440 (W5043, W7065, W7066);
nor G6441 (W5044, W7067, W7068);
nor G6442 (W5045, W7069, W7070);
nor G6443 (W5046, W7071, W7072);
nor G6444 (W5047, W7073, W7074);
nor G6445 (W5048, W7075, W7076);
nor G6446 (W5049, W7077, W7078);
nor G6447 (W5050, W7079, W7080);
nor G6448 (W5051, W7081, W7082);
nor G6449 (W5052, W7083, W7084);
nor G6450 (W5053, W7085, W7086);
nor G6451 (W5054, W7087, W7088);
nor G6452 (W5055, W7089, W7090);
nor G6453 (W5056, W7091, W7092);
nor G6454 (W5057, W7093, W7094);
nor G6455 (W5058, W7095, W7096);
nor G6456 (W5059, W7097, W7098);
nor G6457 (W5060, W7099, W7100);
nor G6458 (W5061, W7101, W7102);
nor G6459 (W5062, W7103, W7104);
nor G6460 (W5063, W7105, W7106);
nor G6461 (W5064, W7107, W7108);
nor G6462 (W5065, W7109, W7110);
nor G6463 (W5066, W7111, W7112);
nor G6464 (W5067, W7113, W7114);
nor G6465 (W5068, W7115, W7116);
nor G6466 (W5069, W7117, W7118);
nor G6467 (W5070, W7119, W7120);
nor G6468 (W5071, W7121, W7122);
nor G6469 (W5072, W7123, W7124);
nor G6470 (W5073, W7125, W7126);
nor G6471 (W5074, W7127, W7128);
nor G6472 (W5075, W7129, W7130);
nor G6473 (W5076, W7131, W7132);
nor G6474 (W5077, W7133, W7134);
nand G6475 (W5078, W5079, W7135);
not G6476 (W5079, W7136);
nor G6477 (W5080, W7137, W7138);
nor G6478 (W5081, W7139, W7140);
nor G6479 (W5082, W7141, W7142);
nor G6480 (W5083, W7143, W7144);
nor G6481 (W5084, W7145, W7146);
nor G6482 (W5085, W7147, W7148);
nor G6483 (W5086, W7149, W7150);
nor G6484 (W5087, W7151, W7152);
nor G6485 (W5088, W7153, W7154);
nor G6486 (W5089, W7155, W7156);
nor G6487 (W5090, W7157, W7158);
nor G6488 (W5091, W7159, W7160);
nor G6489 (W5092, W7161, W7162);
nor G6490 (W5093, W7163, W7164);
nor G6491 (W5094, W7165, W7166);
nor G6492 (W5095, W7167, W7168);
nor G6493 (W5096, W7169, W7170);
nor G6494 (W5097, W7171, W7172);
nor G6495 (W5098, W7173, W7174);
nor G6496 (W5099, W7175, W7176);
nor G6497 (W5100, W7177, W7178);
nor G6498 (W5101, W7179, W7180);
nor G6499 (W5102, W7181, W7182);
nor G6500 (W5103, W7183, W7184);
nor G6501 (W5104, W7185, W7186);
nor G6502 (W5105, W7187, W7188);
nor G6503 (W5106, W7189, W7190);
nor G6504 (W5107, W7191, W7192);
nor G6505 (W5108, W7193, W7194);
nor G6506 (W5109, W7195, W7196);
not G6507 (W5110, W7197);
not G6508 (W5111, W7198);
not G6509 (W5112, W7199);
not G6510 (W5113, W7200);
not G6511 (W5114, W7201);
not G6512 (W5115, W7202);
not G6513 (W5116, W7203);
not G6514 (W5117, W7204);
not G6515 (W5118, W7205);
not G6516 (W5119, W7206);
not G6517 (W5120, W7207);
not G6518 (W5121, W7208);
not G6519 (W5122, W7209);
not G6520 (W5123, W7210);
not G6521 (W5124, W7211);
not G6522 (W5125, W7212);
not G6523 (W5126, W7213);
nor G6524 (W5127, W7214, W7215);
nor G6525 (W5128, W7216, W7217);
nor G6526 (W5129, W7218, W7219);
nor G6527 (W5130, W7220, W7221);
nor G6528 (W5131, W7222, W7223);
nor G6529 (W5132, W7224, W7225);
nor G6530 (W5133, W7226, W7227);
nor G6531 (W5134, W7228, W7229);
nor G6532 (W5135, W7230, W7231);
nor G6533 (W5136, W7232, W7233);
nor G6534 (W5137, W7234, W7235);
nor G6535 (W5138, W7236, W7237);
nor G6536 (W5139, W7238, W7239);
nor G6537 (W5140, W7240, W7241);
nor G6538 (W5141, W7242, W7243);
nor G6539 (W5142, W7244, W7245);
nor G6540 (W5143, W7246, W7247);
nor G6541 (W5144, W7248, W7249);
nor G6542 (W5145, W7250, W7251);
nor G6543 (W5146, W7252, W7253);
nor G6544 (W5147, W7254, W7255);
nor G6545 (W5148, W7256, W7257);
nor G6546 (W5149, W7258, W7259);
nor G6547 (W5150, W7260, W7261);
nor G6548 (W5151, W7262, W7263);
nor G6549 (W5152, W7264, W7265);
nor G6550 (W5153, W7266, W7267);
nor G6551 (W5154, W7268, W7269);
nor G6552 (W5155, W7270, W7271);
nor G6553 (W5156, W7272, W7273);
nor G6554 (W5157, W7274, W7275);
nor G6555 (W5158, W7276, W7275);
nor G6556 (W5159, W7277, W7275);
nor G6557 (W5160, W7278, W7275);
nor G6558 (W5161, W7279, W7275);
nor G6559 (W5162, W7280, W7275);
nor G6560 (W5163, W7281, W7275);
nor G6561 (W5164, W7282, W7275);
nor G6562 (W5165, W7283, W7275);
nor G6563 (W5166, W7284, W7275);
not G6564 (W5167, W7285);
nor G6565 (W5168, W7286, W7287);
nor G6566 (W5169, W7288, W7289);
nor G6567 (W5170, W7290, W7291);
nor G6568 (W5171, W7292, W7293);
nor G6569 (W5172, W7294, W7295);
nor G6570 (W5173, W7296, W7297);
nor G6571 (W5174, W7298, W7299);
nor G6572 (W5175, W7300, W7301);
nor G6573 (W5176, W7302, W7303);
nor G6574 (W5177, W7304, W7305);
nor G6575 (W5178, W7306, W7307);
nor G6576 (W5179, W7308, W7309);
not G6577 (W5180, W7310);
not G6578 (W5181, W7311);
not G6579 (W5182, W7312);
not G6580 (W5183, W7313);
not G6581 (W5184, W7314);
not G6582 (W5185, W7315);
not G6583 (W5186, W7316);
not G6584 (W5187, W7317);
not G6585 (W5188, W7318);
nor G6586 (W5189, W7319, W7320);
nor G6587 (W5190, W7321, W7322);
nor G6588 (W5191, W7323, W7324);
nor G6589 (W5192, W7325, W7326);
nor G6590 (W5193, W7327, W7328);
nor G6591 (W5194, W7329, W7330);
nor G6592 (W5195, W7331, W7332);
nor G6593 (W5196, W7333, W7334);
nor G6594 (W5197, W7335, W7336);
nor G6595 (W5198, W7337, W7338);
nor G6596 (W5199, W7339, W7340);
nor G6597 (W5200, W7341, W7342);
nor G6598 (W5201, W7343, W7344);
nor G6599 (W5202, W7345, W7346);
nor G6600 (W5203, W7347, W7348);
nor G6601 (W5204, W7349, W7350);
nor G6602 (W5205, W7351, W7352);
nor G6603 (W5206, W7353, W7354);
nor G6604 (W5207, W7355, W7356);
nor G6605 (W5208, W7357, W7358);
nor G6606 (W5209, W7359, W7360);
nor G6607 (W5210, W7361, W7362);
nor G6608 (W5211, W7363, W7364);
nor G6609 (W5212, W7365, W7366);
nor G6610 (W5213, W7367, W7368);
nor G6611 (W5214, W7369, W7370);
nor G6612 (W5215, W7371, W7372);
nor G6613 (W5216, W7373, W7374);
nor G6614 (W5217, W7375, W7376);
nor G6615 (W5218, W7377, W7378);
nor G6616 (W5219, W7379, W7380);
nor G6617 (W5220, W7381, W7382);
nor G6618 (W5221, W7383, W7384);
nor G6619 (W5222, W7385, W7386);
nor G6620 (W5223, W7387, W7388);
nor G6621 (W5224, W7389, W7390);
nor G6622 (W5225, W7391, W7392);
nor G6623 (W5226, W7393, W7394);
nor G6624 (W5227, W7395, W7396);
nor G6625 (W5228, W7397, W7398);
nor G6626 (W5229, W7399, W7400);
nor G6627 (W5230, W7401, W7402);
nor G6628 (W5231, W7403, W7404);
nor G6629 (W5232, W7405, W7404);
nor G6630 (W5233, W7406, W7404);
nor G6631 (W5234, W7407, W7404);
nor G6632 (W5235, W7408, W7404);
nor G6633 (W5236, W7409, W7404);
nor G6634 (W5237, W7410, W7404);
nor G6635 (W5238, W7411, W7404);
nor G6636 (W5239, W7412, W7404);
nor G6637 (W5240, W7413, W7404);
nor G6638 (W5241, W7414, W7415);
nor G6639 (W5242, W7416, W7417);
nor G6640 (W5243, W7418, W7419);
nor G6641 (W5244, W7420, W7421);
nor G6642 (W5245, W7422, W7423);
nor G6643 (W5246, W7424, W7425);
nor G6644 (W5247, W7426, W7427);
nor G6645 (W5248, W7428, W7429);
nor G6646 (W5249, W7430, W7431);
not G6647 (W5250, W7432);
not G6648 (W5251, W7433);
not G6649 (W5252, W7434);
not G6650 (W5253, W7435);
nor G6651 (W5254, W7436, W7437);
nor G6652 (W5255, W7438, W7439);
nor G6653 (W5256, W7440, W7441);
nor G6654 (W5257, W7442, W7443);
nor G6655 (W5258, W7444, W7445);
nor G6656 (W5259, W7446, W7447);
nor G6657 (W5260, W7448, W7449);
nor G6658 (W5261, W7450, W7451);
nor G6659 (W5262, W7452, W7453);
nor G6660 (W5263, W7454, W7455);
not G6661 (W5264, W7456);
nor G6662 (W5265, W7457, W7458);
not G6663 (W5266, W7459);
nor G6664 (W5267, W7460, W7461);
not G6665 (W5268, W7462);
nor G6666 (W5269, W7463, W7464);
not G6667 (W5270, W7465);
nor G6668 (W5271, W7466, W7467);
nor G6669 (W5272, W7468, W7469);
nor G6670 (W5273, W7470, W7471);
not G6671 (W5274, W7472);
nor G6672 (W5275, W7473, W7474);
nor G6673 (W5276, W7475, W7476);
nor G6674 (W5277, W7477, W7478);
not G6675 (W5278, W7479);
nor G6676 (W5279, W7480, W7481);
not G6677 (W5280, W7482);
nor G6678 (W5281, W7483, W7484);
nor G6679 (W5282, W7485, W7486);
not G6680 (W5283, W7487);
not G6681 (W5284, W7488);
nor G6682 (W5285, W7489, W7490);
nor G6683 (W5286, W7491, W7492);
nor G6684 (W5287, W7493, W7494);
nor G6685 (W5288, W7495, W7496, W7497);
nor G6686 (W5289, W7498, W7499, W7500);
nor G6687 (W5290, W7501, W7502);
nor G6688 (W5291, W7503, W7504);
nor G6689 (W5292, W7505, W7506);
nor G6690 (W5293, W7507, W7508);
nor G6691 (W5294, W7509, W7510);
nor G6692 (W5295, W7511, W7512);
nor G6693 (W5296, W7513, W7514);
nor G6694 (W5297, W7515, W7516);
not G6695 (W5298, W7517);
not G6696 (W5299, W7518);
not G6697 (W5300, W7519);
not G6698 (W5301, W7520);
not G6699 (W5302, W7521);
not G6700 (W5303, W7522);
not G6701 (W5304, W7523);
not G6702 (W5305, W7524);
not G6703 (W5306, W7525);
not G6704 (W5307, W7526);
nor G6705 (W5308, W7527, W7528);
nor G6706 (W5309, W7529, W7530);
nor G6707 (W5310, W7531, W7532);
nor G6708 (W5311, W7533, W7534);
nor G6709 (W5312, W7535, W7536);
nor G6710 (W5313, W7537, W7538);
nor G6711 (W5314, W7539, W7540);
nor G6712 (W5315, W7541, W7542);
nor G6713 (W5316, W7543, W7544);
nor G6714 (W5317, W7545, W7546);
nor G6715 (W5318, W7547, W7548);
nor G6716 (W5319, W7549, W7550);
nor G6717 (W5320, W7551, W7552);
nor G6718 (W5321, W7553, W7554);
nor G6719 (W5322, W7555, W7556);
nor G6720 (W5323, W7557, W7558);
nor G6721 (W5324, W7559, W7560);
nor G6722 (W5325, W7561, W7562);
nor G6723 (W5326, W7563, W7564);
nor G6724 (W5327, W7565, W7566);
nor G6725 (W5328, W7567, W7568);
nor G6726 (W5329, W7569, W7570);
nor G6727 (W5330, W7571, W7572);
nor G6728 (W5331, W7573, W7574);
nor G6729 (W5332, W7575, W7576);
nor G6730 (W5333, W7577, W7578);
nor G6731 (W5334, W7579, W7580);
nor G6732 (W5335, W7581, W7582);
nor G6733 (W5336, W7583, W7584);
nor G6734 (W5337, W7585, W7586);
nor G6735 (W5338, W7587, W7588);
nor G6736 (W5339, W7589, W7590);
nor G6737 (W5340, W7591, W7592);
nor G6738 (W5341, W7593, W7594);
nor G6739 (W5342, W7595, W7596);
nor G6740 (W5343, W7597, W7598);
nor G6741 (W5344, W7599, W7600);
nor G6742 (W5345, W7601, W7602);
nor G6743 (W5346, W7603, W7604);
nor G6744 (W5347, W7605, W7606);
nor G6745 (W5348, W7607, W7608);
nor G6746 (W5349, W7609, W7610);
nor G6747 (W5350, W7611, W7612);
nor G6748 (W5351, W7613, W7614);
nor G6749 (W5352, W7615, W7616);
nand G6750 (W5353, W5354, W7617);
not G6751 (W5354, W7618);
nor G6752 (W5355, W7619, W7620);
nor G6753 (W5356, W7621, W7622);
nor G6754 (W5357, W7623, W7624);
nor G6755 (W5358, W7625, W7626);
nor G6756 (W5359, W7627, W7628);
nor G6757 (W5360, W7629, W7630);
nor G6758 (W5361, W7631, W7632);
nor G6759 (W5362, W7633, W7634);
nor G6760 (W5363, W7635, W7636);
nor G6761 (W5364, W7637, W7638);
nor G6762 (W5365, W7639, W7640);
nor G6763 (W5366, W7641, W7642);
nor G6764 (W5367, W7643, W7644);
nor G6765 (W5368, W7645, W7646);
nor G6766 (W5369, W7647, W7648);
nor G6767 (W5370, W7649, W7650);
nor G6768 (W5371, W7651, W7652);
nor G6769 (W5372, W7653, W7654);
nor G6770 (W5373, W7655, W7656);
nor G6771 (W5374, W7657, W7658);
nor G6772 (W5375, W7659, W7660);
nor G6773 (W5376, W7661, W7662);
nor G6774 (W5377, W7663, W7664);
nor G6775 (W5378, W7665, W7666);
nor G6776 (W5379, W7667, W7668);
nor G6777 (W5380, W7669, W7670);
nor G6778 (W5381, W7671, W7672);
nor G6779 (W5382, W7673, W7674);
nor G6780 (W5383, W7675, W7676);
nor G6781 (W5384, W7677, W7678);
not G6782 (W5385, W7679);
not G6783 (W5386, W7680);
not G6784 (W5387, W7681);
not G6785 (W5388, W7682);
not G6786 (W5389, W7683);
not G6787 (W5390, W7684);
not G6788 (W5391, W7685);
not G6789 (W5392, W7686);
not G6790 (W5393, W7687);
not G6791 (W5394, W7688);
not G6792 (W5395, W7689);
not G6793 (W5396, W7690);
not G6794 (W5397, W7691);
not G6795 (W5398, W7692);
not G6796 (W5399, W7693);
not G6797 (W5400, W7694);
not G6798 (W5401, W7695);
nor G6799 (W5402, W7696, W7697);
nor G6800 (W5403, W7698, W7699);
nor G6801 (W5404, W7700, W7701);
nor G6802 (W5405, W7702, W7703);
nor G6803 (W5406, W7704, W7705);
nor G6804 (W5407, W7706, W7707);
nor G6805 (W5408, W7708, W7709);
nor G6806 (W5409, W7710, W7711);
nor G6807 (W5410, W7712, W7713);
nor G6808 (W5411, W7714, W7715);
nor G6809 (W5412, W7716, W7717);
nor G6810 (W5413, W7718, W7719);
nor G6811 (W5414, W7720, W7721);
nor G6812 (W5415, W7722, W7723);
nor G6813 (W5416, W7724, W7725);
nor G6814 (W5417, W7726, W7727);
nor G6815 (W5418, W7728, W7729);
nor G6816 (W5419, W7730, W7731);
nor G6817 (W5420, W7732, W7733);
nor G6818 (W5421, W7734, W7735);
nor G6819 (W5422, W7736, W7737);
nor G6820 (W5423, W7738, W7739);
nor G6821 (W5424, W7740, W7741);
nor G6822 (W5425, W7742, W7743);
nor G6823 (W5426, W7744, W7745);
nor G6824 (W5427, W7746, W7747);
nor G6825 (W5428, W7748, W7749);
nor G6826 (W5429, W7750, W7751);
nor G6827 (W5430, W7752, W7753);
nor G6828 (W5431, W7754, W7755);
nor G6829 (W5432, W7756, W7757);
nor G6830 (W5433, W7758, W7757);
nor G6831 (W5434, W7759, W7757);
nor G6832 (W5435, W7760, W7757);
nor G6833 (W5436, W7761, W7757);
nor G6834 (W5437, W7762, W7757);
nor G6835 (W5438, W7763, W7757);
nor G6836 (W5439, W7764, W7757);
nor G6837 (W5440, W7765, W7757);
nor G6838 (W5441, W7766, W7757);
not G6839 (W5442, W7767);
nor G6840 (W5443, W7768, W7769);
nor G6841 (W5444, W7770, W7771);
nor G6842 (W5445, W7772, W7773);
nor G6843 (W5446, W7774, W7775);
nor G6844 (W5447, W7776, W7777);
nor G6845 (W5448, W7778, W7779);
nor G6846 (W5449, W7780, W7781);
nor G6847 (W5450, W7782, W7783);
nor G6848 (W5451, W7784, W7785);
nor G6849 (W5452, W7786, W7787);
nor G6850 (W5453, W7788, W7789);
nor G6851 (W5454, W7790, W7791);
not G6852 (W5455, W7792);
not G6853 (W5456, W7793);
nor G6854 (W5457, W7794, W7795);
nor G6855 (W5458, W7796, W7797);
nor G6856 (W5459, W7798, W7799);
nor G6857 (W5460, W7800, W7801);
not G6858 (W5461, W7802);
not G6859 (W5462, W7803);
not G6860 (W5463, W5462);
not G6861 (W5464, W7804);
not G6862 (W5465, W7805);
not G6863 (W5466, W5465);
not G6864 (W5467, W7806);
not G6865 (W5468, I223);
nor G6866 (W5469, W7807, W7808);
not G6867 (W5470, I224);
nor G6868 (W5471, W7809, W7810);
not G6869 (W5472, I225);
nor G6870 (W5473, W7811, W7812);
not G6871 (W5474, I226);
nor G6872 (W5475, W7813, W7814);
not G6873 (W5476, I227);
nor G6874 (W5477, W7815, W7816);
nor G6875 (W5478, W7817, W7818);
not G6876 (W5479, I228);
not G6877 (W5480, I229);
nor G6878 (W5481, W7819, W7820);
not G6879 (W5482, I230);
nor G6880 (W5483, W7821, W7822);
not G6881 (W5484, W7823);
not G6882 (W5485, I231);
nor G6883 (W5486, W7824, W7825);
not G6884 (W5487, I232);
nor G6885 (W5488, W7826, W7827);
not G6886 (W5489, I233);
nor G6887 (W5490, W7828, W7829);
not G6888 (W5491, I234);
nor G6889 (W5492, W7830, W7831);
not G6890 (W5493, I235);
nor G6891 (W5494, W7832, W7833);
not G6892 (W5495, I236);
nor G6893 (W5496, W7834, W7835);
not G6894 (W5497, I237);
nor G6895 (W5498, W7836, W7837);
not G6896 (W5499, I238);
nor G6897 (W5500, W7838, W7839);
not G6898 (W5501, W7840);
not G6899 (W5502, I239);
nor G6900 (W5503, W7841, W7842);
not G6901 (W5504, I240);
nor G6902 (W5505, W7843, W7844);
not G6903 (W5506, I241);
nor G6904 (W5507, W7845, W7846);
not G6905 (W5508, I242);
nor G6906 (W5509, W7847, W7848);
not G6907 (W5510, I243);
nor G6908 (W5511, W7849, W7850);
not G6909 (W5512, I244);
nor G6910 (W5513, W7851, W7852);
not G6911 (W5514, I245);
nor G6912 (W5515, W7853, W7854);
not G6913 (W5516, I246);
nor G6914 (W5517, W7855, W7856);
not G6915 (W5518, W7857);
nor G6916 (W5519, W7858, W7859);
not G6917 (W5520, I247);
not G6918 (W5521, I248);
nor G6919 (W5522, W7860, W7861);
not G6920 (W5523, I249);
nor G6921 (W5524, W7862, W7863);
not G6922 (W5525, I250);
nor G6923 (W5526, W7864, W7865);
nor G6924 (W5527, W7866, W7867);
not G6925 (W5528, I251);
nor G6926 (W5529, W7868, W7869);
not G6927 (W5530, I252);
not G6928 (W5531, I253);
nor G6929 (W5532, W7870, W7871);
not G6930 (W5533, I254);
nor G6931 (W5534, W7872, W7873);
nand G6932 (W5535, W7874, W7875);
nand G6933 (W5536, W7876, W7877);
nand G6934 (W5537, I255, W7878);
not G6935 (W5538, W7879);
not G6936 (W5539, W7880);
not G6937 (W5540, W7881);
not G6938 (W5541, W7882);
nor G6939 (W5542, W7883, W7884);
nor G6940 (W5543, W7885, W7884);
nor G6941 (W5544, W7886, W7884);
nand G6942 (W5545, W7887, W7888);
nor G6943 (W5546, W7889, W7890);
nor G6944 (W5547, W7891, W7890);
nor G6945 (W5548, W7892, W7890);
nor G6946 (W5549, W7893, W7890);
nor G6947 (W5550, W7894, W7890);
nor G6948 (W5551, W7895, W7890);
nand G6949 (W5552, W7896, W7897);
nor G6950 (W5553, W7898, W7899);
not G6951 (W5554, W7900);
not G6952 (W5555, W7901);
not G6953 (W5556, W7902);
not G6954 (W5557, W7903);
not G6955 (W5558, W7904);
not G6956 (W5559, W7905);
not G6957 (W5560, W7906);
not G6958 (W5561, W7907);
not G6959 (W5562, W7908);
not G6960 (W5563, W7909);
not G6961 (W5564, W7910);
not G6962 (W5565, W7911);
nand G6963 (W5566, W7912, W7913);
nor G6964 (W5567, W7914, W7898);
not G6965 (W5568, W7915);
not G6966 (W5569, W7916);
nand G6967 (W5570, W7917, W7918);
nand G6968 (W5571, W7919, W7920);
nand G6969 (W5572, W7921, W7920);
nand G6970 (W5573, W7922, W7923);
nand G6971 (W5574, W7924, W7925);
nand G6972 (W5575, W7921, W7925);
and G6973 (W5576, W7926, W7927);
and G6974 (W5577, W7928, W7929);
and G6975 (W5578, W7930, W7931);
and G6976 (W5579, W7932, W7933);
and G6977 (W5580, W7934, W7935);
and G6978 (W5581, W7936, W7937);
and G6979 (W5582, W7938, W7939);
and G6980 (W5583, W7940, W7941);
and G6981 (W5584, W7942, W7943);
and G6982 (W5585, W7944, W7945);
and G6983 (W5586, W7946, W7947);
and G6984 (W5587, W7948, W7949);
and G6985 (W5588, W7950, W7951);
and G6986 (W5589, W7952, W7953);
and G6987 (W5590, W7954, W7955);
and G6988 (W5591, W7956, W7957);
and G6989 (W5592, W7958, W7959);
and G6990 (W5593, W7960, W7961);
and G6991 (W5594, W7962, W7963);
and G6992 (W5595, W7964, W7965);
and G6993 (W5596, W7966, W7967);
and G6994 (W5597, W7968, W7969);
and G6995 (W5598, W7970, W7971);
and G6996 (W5599, W7972, W7973);
and G6997 (W5600, W7974, W7975);
and G6998 (W5601, W7976, W7977);
and G6999 (W5602, W7978, W7979);
and G7000 (W5603, W7980, W7981);
and G7001 (W5604, W7982, W7983);
and G7002 (W5605, W7984, W7985);
and G7003 (W5606, W7986, W7987);
and G7004 (W5607, W7988, W7989);
and G7005 (W5608, W7990, W7991);
and G7006 (W5609, W7992, W7993);
and G7007 (W5610, W7994, W7995);
and G7008 (W5611, W7996, W7997);
not G7009 (W5612, W7998);
or G7010 (W5613, I256, W7999);
and G7011 (W5614, W8000, W8001);
and G7012 (W5615, W8002, W8003);
and G7013 (W5616, W8004, W8005);
and G7014 (W5617, W8006, W8007);
and G7015 (W5618, W8008, W8009);
and G7016 (W5619, W8010, W8011);
and G7017 (W5620, W8012, W8013);
and G7018 (W5621, W8014, W8015);
and G7019 (W5622, W8016, W8017);
and G7020 (W5623, W8018, W8019);
and G7021 (W5624, W8020, W8021);
and G7022 (W5625, W8018, W8022);
and G7023 (W5626, W8023, W8024);
and G7024 (W5627, W8018, W8025);
and G7025 (W5628, W8026, W8027);
and G7026 (W5629, W8028, W8029);
and G7027 (W5630, W8030, W8031);
and G7028 (W5631, W8028, W8032);
and G7029 (W5632, W8033, W8034);
and G7030 (W5633, W8028, W8035);
and G7031 (W5634, W8036, W8037);
and G7032 (W5635, W8038, W8039);
and G7033 (W5636, W8040, W8041);
and G7034 (W5637, W8038, W8042);
and G7035 (W5638, W8043, W8044);
and G7036 (W5639, W8038, W8045);
and G7037 (W5640, W8046, W8047);
and G7038 (W5641, W8048, W8049);
and G7039 (W5642, W8050, W8051);
and G7040 (W5643, W8048, W8052);
and G7041 (W5644, W8053, W8054);
and G7042 (W5645, W8048, W8055);
and G7043 (W5646, W8056, W8057);
and G7044 (W5647, W8058, W8059);
and G7045 (W5648, W8060, W8061);
and G7046 (W5649, W8058, W8062);
and G7047 (W5650, W8063, W8064);
and G7048 (W5651, W8058, W8065);
and G7049 (W5652, W8066, W8067);
and G7050 (W5653, W8068, W8069);
and G7051 (W5654, W8070, W8071);
and G7052 (W5655, W8068, W8072);
and G7053 (W5656, W8073, W8074);
and G7054 (W5657, W8068, W8075);
and G7055 (W5658, W8076, W8077);
and G7056 (W5659, W8078, W8079);
and G7057 (W5660, W8080, W8081);
and G7058 (W5661, W8078, W8082);
and G7059 (W5662, W8083, W8084);
and G7060 (W5663, W8078, W8085);
and G7061 (W5664, W8086, W8087);
and G7062 (W5665, W8088, W8089);
and G7063 (W5666, W8090, W8091);
and G7064 (W5667, W8088, W8092);
and G7065 (W5668, W8093, W8094);
and G7066 (W5669, W8088, W8095);
and G7067 (W5670, W8096, W8097);
and G7068 (W5671, W8098, W8099);
and G7069 (W5672, W8100, W8101);
and G7070 (W5673, W8098, W8102);
and G7071 (W5674, W8103, W8104);
and G7072 (W5675, W8098, W8105);
and G7073 (W5676, W8106, W8107);
and G7074 (W5677, W8108, W8109);
and G7075 (W5678, W8110, W8111);
and G7076 (W5679, W8108, W8112);
and G7077 (W5680, W8113, W8114);
and G7078 (W5681, W8108, W8115);
and G7079 (W5682, W8116, W8117);
and G7080 (W5683, W8118, W8119);
and G7081 (W5684, W8120, W8121);
and G7082 (W5685, W8118, W8122);
and G7083 (W5686, W8123, W8124);
and G7084 (W5687, W8118, W8125);
and G7085 (W5688, W8126, W8127);
and G7086 (W5689, W8128, W8129);
and G7087 (W5690, W8130, W8131);
and G7088 (W5691, W8128, W8132);
and G7089 (W5692, W8133, W8134);
and G7090 (W5693, W8128, W8135);
and G7091 (W5694, W8136, W8137);
and G7092 (W5695, W8138, W8139);
and G7093 (W5696, W8140, W8141);
and G7094 (W5697, W8138, W8142);
and G7095 (W5698, W8143, W8144);
and G7096 (W5699, W8138, W8145);
and G7097 (W5700, W8146, W8147);
and G7098 (W5701, W8148, W8149);
and G7099 (W5702, W8150, W8151);
and G7100 (W5703, W8148, W8152);
and G7101 (W5704, W8153, W8154);
and G7102 (W5705, W8148, W8155);
and G7103 (W5706, W8156, W8157);
and G7104 (W5707, W8158, W8159);
and G7105 (W5708, W8160, W8161);
and G7106 (W5709, W8158, W8162);
and G7107 (W5710, W8163, W8164);
and G7108 (W5711, W8158, W8165);
and G7109 (W5712, W8166, W8167);
and G7110 (W5713, W8168, W8169);
and G7111 (W5714, W8170, W8171);
and G7112 (W5715, W8168, W8172);
and G7113 (W5716, W8173, W8174);
and G7114 (W5717, W8168, W8175);
nor G7115 (W5718, W8176, W8177);
not G7116 (W5719, W5723);
nor G7117 (W5720, W8178, W8179);
nor G7118 (W5721, W8180, W8181);
nor G7119 (W5722, W8182, W8183);
nor G7120 (W5723, W5847, W8184);
and G7121 (W5724, W8185, W8186);
and G7122 (W5725, W8187, W8188);
and G7123 (W5726, W8189, W8190);
and G7124 (W5727, W8191, W8192);
and G7125 (W5728, W8193, W8194);
and G7126 (W5729, W8195, W8196);
and G7127 (W5730, W8197, W8198);
and G7128 (W5731, W8199, W8200);
and G7129 (W5732, W8201, W8202);
and G7130 (W5733, W8203, W8204);
and G7131 (W5734, W8205, W8206);
and G7132 (W5735, W8207, W8208);
and G7133 (W5736, W8209, W8210);
and G7134 (W5737, W8211, W8212);
and G7135 (W5738, W8213, W8214);
and G7136 (W5739, W8215, W8216);
and G7137 (W5740, W8201, W8217);
and G7138 (W5741, W8218, W8219);
and G7139 (W5742, W8201, W8220);
and G7140 (W5743, W8221, W8222);
and G7141 (W5744, W8205, W8223);
and G7142 (W5745, W8224, W8225);
and G7143 (W5746, W8205, W8226);
and G7144 (W5747, W8227, W8228);
and G7145 (W5748, W8209, W8229);
and G7146 (W5749, W8230, W8231);
and G7147 (W5750, W8209, W8232);
and G7148 (W5751, W8233, W8234);
and G7149 (W5752, W8213, W8235);
and G7150 (W5753, W8236, W8237);
and G7151 (W5754, W8213, W8238);
and G7152 (W5755, W8239, W8240);
and G7153 (W5756, W8241, W8242);
and G7154 (W5757, W8243, W8244);
and G7155 (W5758, W8245, W8246);
and G7156 (W5759, W8247, W8248);
and G7157 (W5760, W8249, W8250);
and G7158 (W5761, W8251, W8252);
and G7159 (W5762, W8253, W8254);
and G7160 (W5763, W8255, W8256);
and G7161 (W5764, W8257, W8258);
and G7162 (W5765, W8259, W8260);
and G7163 (W5766, W8245, W8261);
and G7164 (W5767, W8262, W8263);
and G7165 (W5768, W8245, W8264);
and G7166 (W5769, W8265, W8266);
and G7167 (W5770, W8249, W8267);
and G7168 (W5771, W8268, W8269);
and G7169 (W5772, W8249, W8270);
and G7170 (W5773, W8271, W8272);
and G7171 (W5774, W8253, W8273);
and G7172 (W5775, W8274, W8275);
and G7173 (W5776, W8253, W8276);
and G7174 (W5777, W8277, W8278);
and G7175 (W5778, W8257, W8279);
and G7176 (W5779, W8280, W8281);
and G7177 (W5780, W8257, W8282);
and G7178 (W5781, W8283, W8284);
and G7179 (W5782, W8285, W8242);
and G7180 (W5783, W8286, W8287);
and G7181 (W5784, W8288, W8289);
and G7182 (W5785, W8290, W8291);
and G7183 (W5786, W8292, W8293);
and G7184 (W5787, W8294, W8295);
and G7185 (W5788, W8296, W8297);
and G7186 (W5789, W8298, W8299);
and G7187 (W5790, W8300, W8301);
and G7188 (W5791, W8302, W8303);
and G7189 (W5792, W8288, W8304);
and G7190 (W5793, W8305, W8306);
and G7191 (W5794, W8288, W8307);
and G7192 (W5795, W8308, W8309);
and G7193 (W5796, W8292, W8310);
and G7194 (W5797, W8311, W8312);
and G7195 (W5798, W8292, W8313);
and G7196 (W5799, W8314, W8315);
and G7197 (W5800, W8296, W8316);
and G7198 (W5801, W8317, W8318);
and G7199 (W5802, W8296, W8319);
and G7200 (W5803, W8320, W8321);
and G7201 (W5804, W8300, W8322);
and G7202 (W5805, W8323, W8324);
and G7203 (W5806, W8300, W8325);
and G7204 (W5807, W8326, W8327);
and G7205 (W5808, W8328, W8242);
and G7206 (W5809, W8329, W8330);
and G7207 (W5810, W8331, W8332);
and G7208 (W5811, W8333, W8334);
and G7209 (W5812, W8335, W8336);
and G7210 (W5813, W8337, W8338);
and G7211 (W5814, W8339, W8340);
and G7212 (W5815, W8341, W8342);
and G7213 (W5816, W8343, W8344);
and G7214 (W5817, W8345, W8346);
and G7215 (W5818, W8331, W8347);
and G7216 (W5819, W8348, W8349);
and G7217 (W5820, W8331, W8350);
and G7218 (W5821, W8351, W8352);
and G7219 (W5822, W8335, W8353);
and G7220 (W5823, W8354, W8355);
and G7221 (W5824, W8335, W8356);
and G7222 (W5825, W8357, W8358);
and G7223 (W5826, W8339, W8359);
and G7224 (W5827, W8360, W8361);
and G7225 (W5828, W8339, W8362);
and G7226 (W5829, W8363, W8364);
and G7227 (W5830, W8343, W8365);
and G7228 (W5831, W8366, W8367);
and G7229 (W5832, W8343, W8368);
and G7230 (W5833, W8369, W8370);
and G7231 (W5834, W8371, W8242);
and G7232 (W5835, W8372, W8373);
nor G7233 (W5836, W8374, W8375);
not G7234 (W5837, W8376);
and G7235 (W5838, W5847, W8377);
and G7236 (W5839, W8378, W8379);
and G7237 (W5840, W8380, W8381);
and G7238 (W5841, W5862, W8382);
nor G7239 (W5842, W8383, W8384);
nor G7240 (W5843, W8385, W8386);
nor G7241 (W5844, W8387, W8388);
nor G7242 (W5845, W8389, W8390);
not G7243 (W5846, I257);
not G7244 (W5847, W5862);
not G7245 (W5848, W8391);
not G7246 (W5849, W8391);
not G7247 (W5850, W8391);
not G7248 (W5851, W8391);
not G7249 (W5852, W8391);
not G7250 (W5853, W8391);
not G7251 (W5854, W8391);
not G7252 (W5855, W8391);
not G7253 (W5856, W8391);
not G7254 (W5857, W8391);
not G7255 (W5858, W8391);
not G7256 (W5859, W8391);
not G7257 (W5860, W8391);
not G7258 (W5861, I258);
not G7259 (W5862, W8392);
not G7260 (W5863, I259);
nor G7261 (W5864, W8393, W8394);
nor G7262 (W5865, W8395, W8396);
nor G7263 (W5866, W8397, W8398);
nor G7264 (W5867, W8399, W8400);
nor G7265 (W5868, W8401, W8402);
nor G7266 (W5869, W8403, W8404, W8405);
nor G7267 (W5870, W8406, W8407);
nor G7268 (W5871, W8408, W8409);
nor G7269 (W5872, W8410, W8411);
and G7270 (W5873, W8412, W8413);
and G7271 (W5874, W8414, W8415);
and G7272 (W5875, W8412, W8416);
and G7273 (W5876, W8417, W8418);
and G7274 (W5877, W8412, W8419);
and G7275 (W5878, W8420, W8421);
and G7276 (W5879, W8422, W8423);
and G7277 (W5880, W8424, W8425);
and G7278 (W5881, W8422, W8426);
and G7279 (W5882, W8427, W8428);
and G7280 (W5883, W8422, W8429);
and G7281 (W5884, W8430, W8431);
and G7282 (W5885, W8432, W8433);
and G7283 (W5886, W8434, W8435);
and G7284 (W5887, W8432, W8436);
and G7285 (W5888, W8437, W8438);
and G7286 (W5889, W8432, W8439);
and G7287 (W5890, W8440, W8441);
and G7288 (W5891, W8442, W8443);
and G7289 (W5892, W8444, W8445);
and G7290 (W5893, W8442, W8446);
and G7291 (W5894, W8447, W8448);
and G7292 (W5895, W8442, W8449);
and G7293 (W5896, W8450, W8451);
and G7294 (W5897, I260, W8452);
and G7295 (W5898, W8453, W8454);
and G7296 (W5899, I260, W8455);
and G7297 (W5900, W8456, W8457);
and G7298 (W5901, I260, W8458);
and G7299 (W5902, W8459, W8460);
and G7300 (W5903, I261, W8461);
and G7301 (W5904, W8462, W8463);
and G7302 (W5905, I261, W8464);
and G7303 (W5906, W8465, W8466);
and G7304 (W5907, I261, W8467);
and G7305 (W5908, W8468, W8469);
and G7306 (W5909, I262, W8470);
and G7307 (W5910, W8471, W8472);
and G7308 (W5911, I262, W8473);
and G7309 (W5912, W8474, W8475);
and G7310 (W5913, I262, W8476);
and G7311 (W5914, W8477, W8478);
and G7312 (W5915, I263, W8479);
and G7313 (W5916, W8480, W8481);
and G7314 (W5917, I263, W8482);
and G7315 (W5918, W8483, W8484);
and G7316 (W5919, I263, W8485);
and G7317 (W5920, W8486, W8487);
and G7318 (W5921, I264, W8488);
and G7319 (W5922, W8489, W8490);
and G7320 (W5923, I264, W8491);
and G7321 (W5924, W8492, W8493);
and G7322 (W5925, I264, W8494);
and G7323 (W5926, W8495, W8496);
and G7324 (W5927, I265, W8497);
and G7325 (W5928, W8498, W8499);
and G7326 (W5929, I265, W8500);
and G7327 (W5930, W8501, W8502);
and G7328 (W5931, I265, W8503);
and G7329 (W5932, W8504, W8505);
and G7330 (W5933, I266, W8506);
and G7331 (W5934, W8507, W8508);
and G7332 (W5935, I266, W8509);
and G7333 (W5936, W8510, W8511);
and G7334 (W5937, I266, W8512);
and G7335 (W5938, W8513, W8514);
and G7336 (W5939, I267, W8515);
and G7337 (W5940, W8516, W8517);
and G7338 (W5941, I267, W8518);
and G7339 (W5942, W8519, W8520);
and G7340 (W5943, I267, W8521);
and G7341 (W5944, W8522, W8523);
and G7342 (W5945, I268, W8524);
and G7343 (W5946, W8525, W8526);
and G7344 (W5947, I268, W8527);
and G7345 (W5948, W8528, W8529);
and G7346 (W5949, I268, W8530);
and G7347 (W5950, W8531, W8532);
and G7348 (W5951, I269, W8533);
and G7349 (W5952, W8534, W8535);
and G7350 (W5953, I269, W8536);
and G7351 (W5954, W8537, W8538);
and G7352 (W5955, I269, W8539);
and G7353 (W5956, W8540, W8541);
nor G7354 (W5957, W8542, W8543);
and G7355 (W5958, W8412, W8544);
nor G7356 (W5959, W8545, W8546);
nor G7357 (W5960, W8547, W8548);
nor G7358 (W5961, W8549, W8550);
nor G7359 (W5962, W8551, W8552);
nor G7360 (W5963, W8553, W8554);
nor G7361 (W5964, W8555, W8556);
nor G7362 (W5965, W8557, W8558);
nor G7363 (W5966, W8559, W8560);
nor G7364 (W5967, W8561, W8562);
and G7365 (W5968, W8563, W8564);
and G7366 (W5969, W8565, W8566);
and G7367 (W5970, W8567, W8568);
and G7368 (W5971, W8569, W8570);
and G7369 (W5972, W8571, W8572);
and G7370 (W5973, W8573, W8574);
and G7371 (W5974, W8575, W8576);
and G7372 (W5975, W8577, W8578);
and G7373 (W5976, W8579, W8580);
and G7374 (W5977, W8581, W8582);
and G7375 (W5978, W8583, W8584);
and G7376 (W5979, W8585, W8586);
and G7377 (W5980, W8587, W8588);
and G7378 (W5981, W8589, W8590);
and G7379 (W5982, W8591, W8592);
and G7380 (W5983, W8589, W8593);
and G7381 (W5984, W8594, W8595);
and G7382 (W5985, W8589, W8596);
nor G7383 (W5986, W8597, W8598, W8599);
nor G7384 (W5987, W8600, W8601, W8602);
nor G7385 (W5988, W8603, W8604, W8605);
nor G7386 (W5989, W8606, W8607, W8608);
and G7387 (W5990, W8609, W8610);
and G7388 (W5991, W8611, W8612);
and G7389 (W5992, W8613, W8614);
and G7390 (W5993, W8611, W8615);
and G7391 (W5994, W8616, W8617);
and G7392 (W5995, W8611, W8618);
and G7393 (W5996, W8619, W8620);
and G7394 (W5997, W8621, W8622);
and G7395 (W5998, W8623, W8624);
and G7396 (W5999, W8621, W8625);
and G7397 (W6000, W8626, W8627);
and G7398 (W6001, W8621, W8628);
and G7399 (W6002, W8629, W8630);
and G7400 (W6003, W8631, W8632);
and G7401 (W6004, W8633, W8634);
and G7402 (W6005, W8635, W8636);
and G7403 (W6006, W8637, W8638);
and G7404 (W6007, W8635, W8639);
and G7405 (W6008, W8640, W8641);
and G7406 (W6009, W8635, W8642);
not G7407 (W6010, I270);
and G7408 (W6011, W8643, W8644);
and G7409 (W6012, W8645, W8646);
not G7410 (W6013, I271);
and G7411 (W6014, W8647, W8648);
and G7412 (W6015, W8645, W8649);
not G7413 (W6016, I272);
and G7414 (W6017, W8650, W8651);
and G7415 (W6018, W8645, W8652);
not G7416 (W6019, W8653);
and G7417 (W6020, W8654, W8655);
and G7418 (W6021, W8656, W8657);
and G7419 (W6022, W8658, W8659);
and G7420 (W6023, W8656, W8660);
and G7421 (W6024, W8661, W8662);
and G7422 (W6025, W8656, W8663);
not G7423 (W6026, W8664);
and G7424 (W6027, W8665, W8666);
and G7425 (W6028, W8667, W8668);
and G7426 (W6029, W8669, W8670);
and G7427 (W6030, W8667, W8671);
and G7428 (W6031, W8672, W8673);
and G7429 (W6032, W8667, W8674);
not G7430 (W6033, I273);
and G7431 (W6034, W8675, W8676);
and G7432 (W6035, W8677, W8678);
not G7433 (W6036, I274);
and G7434 (W6037, W8679, W8680);
and G7435 (W6038, W8677, W8681);
and G7436 (W6039, W8682, W8683);
and G7437 (W6040, W8677, W8684);
not G7438 (W6041, I275);
not G7439 (W6042, W8685);
and G7440 (W6043, W8686, W8687);
and G7441 (W6044, W8688, W8689);
and G7442 (W6045, W8690, W8691);
and G7443 (W6046, W8688, W8692);
and G7444 (W6047, W8693, W8694);
and G7445 (W6048, W8688, W8695);
and G7446 (W6049, W8696, I276);
and G7447 (W6050, W8697, I277);
and G7448 (W6051, W8698, I278);
and G7449 (W6052, W8696, I279);
and G7450 (W6053, W8697, I280);
and G7451 (W6054, W8698, I281);
and G7452 (W6055, W8699, W8700);
and G7453 (W6056, W8701, W8702);
and G7454 (W6057, W8701, W8703);
and G7455 (W6058, I282, W8704);
and G7456 (W6059, W8705, W8706);
and G7457 (W6060, I283, W8707);
and G7458 (W6061, W8708, W8709);
and G7459 (W6062, W8710, W8711);
and G7460 (W6063, W8712, W8713);
and G7461 (W6064, W8714, W8715);
and G7462 (W6065, W8716, W8717);
and G7463 (W6066, W8718, W8719);
and G7464 (W6067, W8720, W8721);
and G7465 (W6068, W8722, W8723);
and G7466 (W6069, W8724, W8725);
and G7467 (W6070, W8726, W8727);
not G7468 (W6071, W8728);
not G7469 (W6072, W8729);
not G7470 (W6073, W8730);
not G7471 (W6074, W8731);
not G7472 (W6075, W8732);
not G7473 (W6076, W8733);
not G7474 (W6077, W8734);
not G7475 (W6078, W8735);
not G7476 (W6079, W8736);
not G7477 (W6080, W8737);
and G7478 (W6081, W8738, W8739);
and G7479 (W6082, W8740, W8741);
and G7480 (W6083, W8738, W8742);
and G7481 (W6084, W8743, W8744);
and G7482 (W6085, W8738, W8745);
and G7483 (W6086, W8746, W8747);
and G7484 (W6087, W8748, W8749);
and G7485 (W6088, W8750, W8751);
and G7486 (W6089, W8752, W8753);
and G7487 (W6090, W8750, W8754);
and G7488 (W6091, W8755, W8756);
and G7489 (W6092, W8750, W8757);
and G7490 (W6093, W8758, W8759);
and G7491 (W6094, W8760, W8761);
and G7492 (W6095, W8762, W8763);
and G7493 (W6096, W8760, W8764);
and G7494 (W6097, W8765, W8766);
and G7495 (W6098, W8760, W8767);
and G7496 (W6099, W8768, W8769);
and G7497 (W6100, W8770, W8771);
and G7498 (W6101, W8772, W8773);
and G7499 (W6102, W8770, W8774);
and G7500 (W6103, W8775, W8776);
and G7501 (W6104, W8770, W8777);
and G7502 (W6105, W8778, W8779);
and G7503 (W6106, W8780, W8781);
and G7504 (W6107, W8782, W8783);
and G7505 (W6108, W8780, W8784);
and G7506 (W6109, W8785, W8786);
and G7507 (W6110, W8780, W8787);
and G7508 (W6111, W8788, W8789);
and G7509 (W6112, W8790, W8791);
and G7510 (W6113, W8792, W8793);
and G7511 (W6114, W8790, W8794);
and G7512 (W6115, W8795, W8796);
and G7513 (W6116, W8790, W8797);
and G7514 (W6117, W8798, W8799);
and G7515 (W6118, W8800, W8801);
and G7516 (W6119, W8802, W8803);
and G7517 (W6120, W8800, W8804);
and G7518 (W6121, W8805, W8806);
and G7519 (W6122, W8800, W8807);
and G7520 (W6123, W8808, W8809);
and G7521 (W6124, W8810, W8811);
and G7522 (W6125, W8812, W8813);
and G7523 (W6126, W8810, W8814);
and G7524 (W6127, W8815, W8816);
and G7525 (W6128, W8810, W8817);
and G7526 (W6129, W8818, W8819);
and G7527 (W6130, W8820, W8821);
and G7528 (W6131, W8822, W8823);
and G7529 (W6132, W8820, W8824);
and G7530 (W6133, W8825, W8826);
and G7531 (W6134, W8820, W8827);
and G7532 (W6135, W8828, W8829);
and G7533 (W6136, W8830, W8831);
and G7534 (W6137, W8832, W8833);
and G7535 (W6138, W8830, W8834);
and G7536 (W6139, W8835, W8836);
and G7537 (W6140, W8830, W8837);
and G7538 (W6141, W8838, W8839);
and G7539 (W6142, W8840, W8841);
and G7540 (W6143, W8842, W8843);
and G7541 (W6144, W8840, W8844);
and G7542 (W6145, W8845, W8846);
and G7543 (W6146, W8840, W8847);
and G7544 (W6147, W8848, W8849);
and G7545 (W6148, W8850, W8851);
and G7546 (W6149, W8852, W8853);
and G7547 (W6150, W8850, W8854);
and G7548 (W6151, W8855, W8856);
and G7549 (W6152, W8850, W8857);
and G7550 (W6153, W8858, W8859);
and G7551 (W6154, W8860, W8861);
and G7552 (W6155, W8862, W8863);
and G7553 (W6156, W8860, W8864);
and G7554 (W6157, W8865, W8866);
and G7555 (W6158, W8860, W8867);
and G7556 (W6159, W8868, W8869);
and G7557 (W6160, W8870, W8871);
and G7558 (W6161, W8872, W8873);
and G7559 (W6162, W8870, W8874);
and G7560 (W6163, W8875, W8876);
and G7561 (W6164, W8870, W8877);
and G7562 (W6165, W8878, W8879);
and G7563 (W6166, W8880, W8881);
and G7564 (W6167, W8878, W8882);
and G7565 (W6168, W8883, W8884);
and G7566 (W6169, W8878, W8885);
and G7567 (W6170, W8886, W8887);
not G7568 (W6171, W8888);
not G7569 (W6172, W8889);
and G7570 (W6173, W8890, W8891);
and G7571 (W6174, W8892, W8893);
and G7572 (W6175, W8894, W8895);
and G7573 (W6176, W8896, W8897);
and G7574 (W6177, W8898, W8899);
and G7575 (W6178, W8900, W8901);
and G7576 (W6179, W8902, W8903);
and G7577 (W6180, W8904, W8905);
and G7578 (W6181, W8890, W8906);
and G7579 (W6182, W8907, W8908);
and G7580 (W6183, W8890, W8909);
and G7581 (W6184, W8910, W8911);
and G7582 (W6185, W8894, W8912);
and G7583 (W6186, W8913, W8914);
and G7584 (W6187, W8894, W8915);
and G7585 (W6188, W8916, W8917);
and G7586 (W6189, W8898, W8918);
and G7587 (W6190, W8919, W8920);
and G7588 (W6191, W8898, W8921);
and G7589 (W6192, W8922, W8923);
and G7590 (W6193, W8902, W8924);
and G7591 (W6194, W8925, W8926);
and G7592 (W6195, W8902, W8927);
and G7593 (W6196, W8928, W8929);
and G7594 (W6197, W8930, W8931);
and G7595 (W6198, W8932, W8933);
and G7596 (W6199, W8934, W8935);
and G7597 (W6200, W8932, W8936);
and G7598 (W6201, W8937, W8938);
and G7599 (W6202, W8932, W8939);
and G7600 (W6203, W8940, W8941);
and G7601 (W6204, W8942, W8943);
and G7602 (W6205, W8940, W8944);
and G7603 (W6206, W8945, W8946);
and G7604 (W6207, W8940, W8947);
and G7605 (W6208, W8948, W8949);
and G7606 (W6209, W8950, W8951);
and G7607 (W6210, W8952, W8953);
and G7608 (W6211, W8954, W8955);
and G7609 (W6212, W8952, W8956);
and G7610 (W6213, W8957, W8958);
and G7611 (W6214, W8952, W8959);
and G7612 (W6215, W8960, W8961);
and G7613 (W6216, W8962, W8963);
and G7614 (W6217, W8964, W8965);
and G7615 (W6218, W8962, W8966);
and G7616 (W6219, W8967, W8968);
and G7617 (W6220, W8962, W8969);
and G7618 (W6221, W8970, W8971);
and G7619 (W6222, W8972, W8973);
and G7620 (W6223, W8974, W8975);
and G7621 (W6224, W8972, W8976);
and G7622 (W6225, W8977, W8978);
and G7623 (W6226, W8972, W8979);
and G7624 (W6227, W8980, W8981);
and G7625 (W6228, W8982, W8983);
and G7626 (W6229, W8980, W8984);
and G7627 (W6230, W8985, W8986);
and G7628 (W6231, W8980, W8987);
and G7629 (W6232, W8988, W8989);
nor G7630 (W6233, W8990, W8991, W8992);
nor G7631 (W6234, W8993, W8994, W8995);
not G7632 (W6235, I284);
not G7633 (W6236, I285);
not G7634 (W6237, I286);
nor G7635 (W6238, W8996, W8997, W8998);
not G7636 (W6239, I287);
not G7637 (W6240, I288);
not G7638 (W6241, I289);
nor G7639 (W6242, W8999, W9000, W9001);
not G7640 (W6243, I290);
not G7641 (W6244, I291);
not G7642 (W6245, I292);
nor G7643 (W6246, W9002, W9003, W9004);
not G7644 (W6247, I293);
not G7645 (W6248, I294);
not G7646 (W6249, I295);
and G7647 (W6250, W9005, W9006);
and G7648 (W6251, W9007, W9008);
and G7649 (W6252, W9009, W9010);
and G7650 (W6253, W9011, W9012);
and G7651 (W6254, W9013, W9014);
and G7652 (W6255, W9015, W9016);
and G7653 (W6256, W9017, W9018);
and G7654 (W6257, W9019, W9020);
and G7655 (W6258, W9021, W9022);
and G7656 (W6259, W9023, W9024);
and G7657 (W6260, W9025, W9026);
and G7658 (W6261, W9027, W9028);
and G7659 (W6262, W9029, W9030);
and G7660 (W6263, W9031, W9032);
and G7661 (W6264, W9033, W9034);
and G7662 (W6265, W9035, W9036);
and G7663 (W6266, W9037, W9038);
and G7664 (W6267, W9039, W9040);
and G7665 (W6268, W9041, W9042);
and G7666 (W6269, W9043, W9044);
and G7667 (W6270, W9005, W9045);
and G7668 (W6271, W9046, W9047);
and G7669 (W6272, W9005, W9048);
and G7670 (W6273, W9049, W9050);
and G7671 (W6274, W9009, W9051);
and G7672 (W6275, W9052, W9053);
and G7673 (W6276, W9009, W9054);
and G7674 (W6277, W9055, W9056);
and G7675 (W6278, W9013, W9057);
and G7676 (W6279, W9058, W9059);
and G7677 (W6280, W9013, W9060);
and G7678 (W6281, W9061, W9062);
and G7679 (W6282, W9017, W9063);
and G7680 (W6283, W9064, W9065);
and G7681 (W6284, W9017, W9066);
and G7682 (W6285, W9067, W9068);
and G7683 (W6286, W9021, W9069);
and G7684 (W6287, W9070, W9071);
and G7685 (W6288, W9021, W9072);
and G7686 (W6289, W9073, W9074);
and G7687 (W6290, W9025, W9075);
and G7688 (W6291, W9076, W9077);
and G7689 (W6292, W9025, W9078);
and G7690 (W6293, W9079, W9080);
and G7691 (W6294, W9029, W9081);
and G7692 (W6295, W9082, W9083);
and G7693 (W6296, W9033, W9084);
and G7694 (W6297, W9085, W9086);
and G7695 (W6298, W9029, W9087);
and G7696 (W6299, W9088, W9089);
and G7697 (W6300, W9037, W9090);
and G7698 (W6301, W9091, W9092);
and G7699 (W6302, W9033, W9093);
and G7700 (W6303, W9094, W9095);
and G7701 (W6304, W9041, W9096);
and G7702 (W6305, W9097, W9098);
and G7703 (W6306, W9037, W9099);
and G7704 (W6307, W9100, W9101);
and G7705 (W6308, W9041, W9102);
and G7706 (W6309, W9103, W9104);
nor G7707 (W6310, W9105, W9106);
and G7708 (W6311, W9107, W9108, W9109);
nor G7709 (W6312, W9110, W9111);
nor G7710 (W6313, W9112, W9113);
nor G7711 (W6314, W9114, W9115);
nor G7712 (W6315, W9116, W9117);
nor G7713 (W6316, W9118, W9119);
nor G7714 (W6317, W9120, W9121);
nor G7715 (W6318, W9122, W9123);
nor G7716 (W6319, W9124, W9125);
nor G7717 (W6320, W9126, W9127);
not G7718 (W6321, I47);
and G7719 (W6322, W9128, W9129);
and G7720 (W6323, W9130, W9131);
and G7721 (W6324, W9128, W9132);
and G7722 (W6325, W9133, W9134);
and G7723 (W6326, W9128, W9135);
and G7724 (W6327, W9136, W9137);
and G7725 (W6328, W9033, W9138);
and G7726 (W6329, W9139, W9140);
and G7727 (W6330, W9033, W9141);
and G7728 (W6331, W9142, W9143);
and G7729 (W6332, W9033, W9144);
and G7730 (W6333, W9145, W9146);
and G7731 (W6334, W9041, W9147);
and G7732 (W6335, W9148, W9149);
and G7733 (W6336, W9041, W9150);
and G7734 (W6337, W9151, W9152);
and G7735 (W6338, W9041, W9153);
and G7736 (W6339, W9154, W9155);
and G7737 (W6340, W9156, W9157);
and G7738 (W6341, W9158, W9159);
and G7739 (W6342, W9156, W9160);
and G7740 (W6343, W9161, W9162);
and G7741 (W6344, W9156, W9163);
and G7742 (W6345, W9164, W9165);
nor G7743 (W6346, W9166, W9167);
nor G7744 (W6347, W9168, W9169);
nor G7745 (W6348, W9170, W9171);
nor G7746 (W6349, W9172, W9173);
nor G7747 (W6350, W9174, W9175);
nor G7748 (W6351, W9176, W9177, W9178);
nor G7749 (W6352, W9179, W9180);
nor G7750 (W6353, W9181, W9182);
nor G7751 (W6354, W9183, W9184);
and G7752 (W6355, W9185, W9186);
and G7753 (W6356, W9187, W9188);
and G7754 (W6357, W9185, W9189);
and G7755 (W6358, W9190, W9191);
and G7756 (W6359, W9185, W9192);
and G7757 (W6360, W9193, W9194);
and G7758 (W6361, W9195, W9196);
and G7759 (W6362, W9197, W9198);
and G7760 (W6363, W9195, W9199);
and G7761 (W6364, W9200, W9201);
and G7762 (W6365, W9195, W9202);
and G7763 (W6366, W9203, W9204);
and G7764 (W6367, W9205, W9206);
and G7765 (W6368, W9207, W9208);
and G7766 (W6369, W9205, W9209);
and G7767 (W6370, W9210, W9211);
and G7768 (W6371, W9205, W9212);
and G7769 (W6372, W9213, W9214);
and G7770 (W6373, W9215, W9216);
and G7771 (W6374, W9217, W9218);
and G7772 (W6375, W9215, W9219);
and G7773 (W6376, W9220, W9221);
and G7774 (W6377, W9215, W9222);
and G7775 (W6378, W9223, W9224);
and G7776 (W6379, I296, W9225);
and G7777 (W6380, W9226, W9227);
and G7778 (W6381, I296, W9228);
and G7779 (W6382, W9229, W9230);
and G7780 (W6383, I296, W9231);
and G7781 (W6384, W9232, W9233);
and G7782 (W6385, I297, W9234);
and G7783 (W6386, W9235, W9236);
and G7784 (W6387, I297, W9237);
and G7785 (W6388, W9238, W9239);
and G7786 (W6389, I297, W9240);
and G7787 (W6390, W9241, W9242);
and G7788 (W6391, I298, W9243);
and G7789 (W6392, W9244, W9245);
and G7790 (W6393, I298, W9246);
and G7791 (W6394, W9247, W9248);
and G7792 (W6395, I298, W9249);
and G7793 (W6396, W9250, W9251);
and G7794 (W6397, I299, W9252);
and G7795 (W6398, W9253, W9254);
and G7796 (W6399, I299, W9255);
and G7797 (W6400, W9256, W9257);
and G7798 (W6401, I299, W9258);
and G7799 (W6402, W9259, W9260);
and G7800 (W6403, I300, W9261);
and G7801 (W6404, W9262, W9263);
and G7802 (W6405, I300, W9264);
and G7803 (W6406, W9265, W9266);
and G7804 (W6407, I300, W9267);
and G7805 (W6408, W9268, W9269);
and G7806 (W6409, I301, W9270);
and G7807 (W6410, W9271, W9272);
and G7808 (W6411, I301, W9273);
and G7809 (W6412, W9274, W9275);
and G7810 (W6413, I301, W9276);
and G7811 (W6414, W9277, W9278);
and G7812 (W6415, I302, W9279);
and G7813 (W6416, W9280, W9281);
and G7814 (W6417, I302, W9282);
and G7815 (W6418, W9283, W9284);
and G7816 (W6419, I302, W9285);
and G7817 (W6420, W9286, W9287);
and G7818 (W6421, I303, W9288);
and G7819 (W6422, W9289, W9290);
and G7820 (W6423, I303, W9291);
and G7821 (W6424, W9292, W9293);
and G7822 (W6425, I303, W9294);
and G7823 (W6426, W9295, W9296);
and G7824 (W6427, I304, W9297);
and G7825 (W6428, W9298, W9299);
and G7826 (W6429, I304, W9300);
and G7827 (W6430, W9301, W9302);
and G7828 (W6431, I304, W9303);
and G7829 (W6432, W9304, W9305);
and G7830 (W6433, I305, W9306);
and G7831 (W6434, W9307, W9308);
and G7832 (W6435, I305, W9309);
and G7833 (W6436, W9310, W9311);
and G7834 (W6437, I305, W9312);
and G7835 (W6438, W9313, W9314);
nor G7836 (W6439, W9315, W9316);
and G7837 (W6440, W9185, W9317);
nor G7838 (W6441, W9318, W9319);
nor G7839 (W6442, W9320, W9321);
nor G7840 (W6443, W9322, W9323);
nor G7841 (W6444, W9324, W9325);
nor G7842 (W6445, W9326, W9327);
nor G7843 (W6446, W9328, W9329);
nor G7844 (W6447, W9330, W9331);
nor G7845 (W6448, W9332, W9333);
nor G7846 (W6449, W9334, W9335);
and G7847 (W6450, W9336, W9337);
and G7848 (W6451, W9338, W9339);
and G7849 (W6452, W9340, W9341);
and G7850 (W6453, W9342, W9343);
and G7851 (W6454, W9344, W9345);
and G7852 (W6455, W9346, W9347);
and G7853 (W6456, W9348, W9349);
and G7854 (W6457, W9350, W9351);
and G7855 (W6458, W9352, W9353);
and G7856 (W6459, W9354, W9355);
and G7857 (W6460, W9356, W9357);
and G7858 (W6461, W9358, W9359);
and G7859 (W6462, W9360, W9361);
and G7860 (W6463, W9362, W9363);
and G7861 (W6464, W9364, W9365);
and G7862 (W6465, W9362, W9366);
and G7863 (W6466, W9367, W9368);
and G7864 (W6467, W9362, W9369);
nor G7865 (W6468, W9370, W9371, W9372);
nor G7866 (W6469, W9373, W9374, W9375);
nor G7867 (W6470, W9376, W9377, W9378);
nor G7868 (W6471, W9379, W9380, W9381);
and G7869 (W6472, W9382, W9383);
and G7870 (W6473, W9384, W9385);
and G7871 (W6474, W9386, W9387);
and G7872 (W6475, W9384, W9388);
and G7873 (W6476, W9389, W9390);
and G7874 (W6477, W9384, W9391);
and G7875 (W6478, W9392, W9393);
and G7876 (W6479, W9394, W9395);
and G7877 (W6480, W9396, W9397);
and G7878 (W6481, W9394, W9398);
and G7879 (W6482, W9399, W9400);
and G7880 (W6483, W9394, W9401);
and G7881 (W6484, W9402, W9403);
and G7882 (W6485, W9404, W9405);
and G7883 (W6486, W9406, W9407);
and G7884 (W6487, W9408, W9409);
and G7885 (W6488, W9410, W9411);
and G7886 (W6489, W9408, W9412);
and G7887 (W6490, W9413, W9414);
and G7888 (W6491, W9408, W9415);
not G7889 (W6492, I306);
and G7890 (W6493, W9416, W9417);
and G7891 (W6494, W9418, W9419);
not G7892 (W6495, I307);
and G7893 (W6496, W9420, W9421);
and G7894 (W6497, W9418, W9422);
not G7895 (W6498, I308);
and G7896 (W6499, W9423, W9424);
and G7897 (W6500, W9418, W9425);
not G7898 (W6501, W9426);
and G7899 (W6502, W9427, W9428);
and G7900 (W6503, W9429, W9430);
and G7901 (W6504, W9431, W9432);
and G7902 (W6505, W9429, W9433);
and G7903 (W6506, W9434, W9435);
and G7904 (W6507, W9429, W9436);
not G7905 (W6508, W9437);
and G7906 (W6509, W9438, W9439);
and G7907 (W6510, W9440, W9441);
and G7908 (W6511, W9442, W9443);
and G7909 (W6512, W9440, W9444);
and G7910 (W6513, W9445, W9446);
and G7911 (W6514, W9440, W9447);
not G7912 (W6515, I309);
and G7913 (W6516, W9448, W9449);
and G7914 (W6517, W9450, W9451);
not G7915 (W6518, I310);
and G7916 (W6519, W9452, W9453);
and G7917 (W6520, W9450, W9454);
and G7918 (W6521, W9455, W9456);
and G7919 (W6522, W9450, W9457);
not G7920 (W6523, I311);
not G7921 (W6524, W9458);
and G7922 (W6525, W9459, W9460);
and G7923 (W6526, W9461, W9462);
and G7924 (W6527, W9463, W9464);
and G7925 (W6528, W9461, W9465);
and G7926 (W6529, W9466, W9467);
and G7927 (W6530, W9461, W9468);
and G7928 (W6531, W9469, I312);
and G7929 (W6532, W9470, I313);
and G7930 (W6533, W9471, I314);
and G7931 (W6534, W9469, I315);
and G7932 (W6535, W9470, I316);
and G7933 (W6536, W9471, I317);
and G7934 (W6537, W9472, W9473);
and G7935 (W6538, W9474, W9475);
and G7936 (W6539, W9474, W9476);
and G7937 (W6540, I318, W9477);
and G7938 (W6541, W9478, W9479);
and G7939 (W6542, I319, W9480);
and G7940 (W6543, W9481, W9482);
and G7941 (W6544, W9483, W9484);
and G7942 (W6545, W9485, W9486);
and G7943 (W6546, W9487, W9488);
and G7944 (W6547, W9489, W9490);
and G7945 (W6548, W9491, W9492);
and G7946 (W6549, W9493, W9494);
and G7947 (W6550, W9495, W9496);
and G7948 (W6551, W9497, W9498);
and G7949 (W6552, W9499, W9500);
not G7950 (W6553, W9501);
not G7951 (W6554, W9502);
not G7952 (W6555, W9503);
not G7953 (W6556, W9504);
not G7954 (W6557, W9505);
not G7955 (W6558, W9506);
not G7956 (W6559, W9507);
not G7957 (W6560, W9508);
not G7958 (W6561, W9509);
not G7959 (W6562, W9510);
and G7960 (W6563, W9511, W9512);
and G7961 (W6564, W9513, W9514);
and G7962 (W6565, W9511, W9515);
and G7963 (W6566, W9516, W9517);
and G7964 (W6567, W9511, W9518);
and G7965 (W6568, W9519, W9520);
and G7966 (W6569, W9521, W9522);
and G7967 (W6570, W9523, W9524);
and G7968 (W6571, W9525, W9526);
and G7969 (W6572, W9523, W9527);
and G7970 (W6573, W9528, W9529);
and G7971 (W6574, W9523, W9530);
and G7972 (W6575, W9531, W9532);
and G7973 (W6576, W9533, W9534);
and G7974 (W6577, W9535, W9536);
and G7975 (W6578, W9533, W9537);
and G7976 (W6579, W9538, W9539);
and G7977 (W6580, W9533, W9540);
and G7978 (W6581, W9541, W9542);
and G7979 (W6582, W9543, W9544);
and G7980 (W6583, W9545, W9546);
and G7981 (W6584, W9543, W9547);
and G7982 (W6585, W9548, W9549);
and G7983 (W6586, W9543, W9550);
and G7984 (W6587, W9551, W9552);
and G7985 (W6588, W9553, W9554);
and G7986 (W6589, W9555, W9556);
and G7987 (W6590, W9553, W9557);
and G7988 (W6591, W9558, W9559);
and G7989 (W6592, W9553, W9560);
and G7990 (W6593, W9561, W9562);
and G7991 (W6594, W9563, W9564);
and G7992 (W6595, W9565, W9566);
and G7993 (W6596, W9563, W9567);
and G7994 (W6597, W9568, W9569);
and G7995 (W6598, W9563, W9570);
and G7996 (W6599, W9571, W9572);
and G7997 (W6600, W9573, W9574);
and G7998 (W6601, W9575, W9576);
and G7999 (W6602, W9573, W9577);
and G8000 (W6603, W9578, W9579);
and G8001 (W6604, W9573, W9580);
and G8002 (W6605, W9581, W9582);
and G8003 (W6606, W9583, W9584);
and G8004 (W6607, W9585, W9586);
and G8005 (W6608, W9583, W9587);
and G8006 (W6609, W9588, W9589);
and G8007 (W6610, W9583, W9590);
and G8008 (W6611, W9591, W9592);
and G8009 (W6612, W9593, W9594);
and G8010 (W6613, W9595, W9596);
and G8011 (W6614, W9593, W9597);
and G8012 (W6615, W9598, W9599);
and G8013 (W6616, W9593, W9600);
and G8014 (W6617, W9601, W9602);
and G8015 (W6618, W9603, W9604);
and G8016 (W6619, W9605, W9606);
and G8017 (W6620, W9603, W9607);
and G8018 (W6621, W9608, W9609);
and G8019 (W6622, W9603, W9610);
and G8020 (W6623, W9611, W9612);
and G8021 (W6624, W9613, W9614);
and G8022 (W6625, W9615, W9616);
and G8023 (W6626, W9613, W9617);
and G8024 (W6627, W9618, W9619);
and G8025 (W6628, W9613, W9620);
and G8026 (W6629, W9621, W9622);
and G8027 (W6630, W9623, W9624);
and G8028 (W6631, W9625, W9626);
and G8029 (W6632, W9623, W9627);
and G8030 (W6633, W9628, W9629);
and G8031 (W6634, W9623, W9630);
and G8032 (W6635, W9631, W9632);
and G8033 (W6636, W9633, W9634);
and G8034 (W6637, W9635, W9636);
and G8035 (W6638, W9633, W9637);
and G8036 (W6639, W9638, W9639);
and G8037 (W6640, W9633, W9640);
and G8038 (W6641, W9641, W9642);
and G8039 (W6642, W9643, W9644);
and G8040 (W6643, W9645, W9646);
and G8041 (W6644, W9643, W9647);
and G8042 (W6645, W9648, W9649);
and G8043 (W6646, W9643, W9650);
and G8044 (W6647, W9651, W9652);
and G8045 (W6648, W9653, W9654);
and G8046 (W6649, W9651, W9655);
and G8047 (W6650, W9656, W9657);
and G8048 (W6651, W9651, W9658);
and G8049 (W6652, W9659, W9660);
not G8050 (W6653, W9661);
not G8051 (W6654, W9662);
and G8052 (W6655, W9663, W9664);
and G8053 (W6656, W9665, W9666);
and G8054 (W6657, W9667, W9668);
and G8055 (W6658, W9669, W9670);
and G8056 (W6659, W9671, W9672);
and G8057 (W6660, W9673, W9674);
and G8058 (W6661, W9675, W9676);
and G8059 (W6662, W9677, W9678);
and G8060 (W6663, W9663, W9679);
and G8061 (W6664, W9680, W9681);
and G8062 (W6665, W9663, W9682);
and G8063 (W6666, W9683, W9684);
and G8064 (W6667, W9667, W9685);
and G8065 (W6668, W9686, W9687);
and G8066 (W6669, W9667, W9688);
and G8067 (W6670, W9689, W9690);
and G8068 (W6671, W9671, W9691);
and G8069 (W6672, W9692, W9693);
and G8070 (W6673, W9671, W9694);
and G8071 (W6674, W9695, W9696);
and G8072 (W6675, W9675, W9697);
and G8073 (W6676, W9698, W9699);
and G8074 (W6677, W9675, W9700);
and G8075 (W6678, W9701, W9702);
and G8076 (W6679, W9703, W9704);
and G8077 (W6680, W9705, W9706);
and G8078 (W6681, W9707, W9708);
and G8079 (W6682, W9705, W9709);
and G8080 (W6683, W9710, W9711);
and G8081 (W6684, W9705, W9712);
and G8082 (W6685, W9713, W9714);
and G8083 (W6686, W9715, W9716);
and G8084 (W6687, W9713, W9717);
and G8085 (W6688, W9718, W9719);
and G8086 (W6689, W9713, W9720);
and G8087 (W6690, W9721, W9722);
and G8088 (W6691, W9723, W9724);
and G8089 (W6692, W9725, W9726);
and G8090 (W6693, W9727, W9728);
and G8091 (W6694, W9725, W9729);
and G8092 (W6695, W9730, W9731);
and G8093 (W6696, W9725, W9732);
and G8094 (W6697, W9733, W9734);
and G8095 (W6698, W9735, W9736);
and G8096 (W6699, W9737, W9738);
and G8097 (W6700, W9735, W9739);
and G8098 (W6701, W9740, W9741);
and G8099 (W6702, W9735, W9742);
and G8100 (W6703, W9743, W9744);
and G8101 (W6704, W9745, W9746);
and G8102 (W6705, W9747, W9748);
and G8103 (W6706, W9745, W9749);
and G8104 (W6707, W9750, W9751);
and G8105 (W6708, W9745, W9752);
and G8106 (W6709, W9753, W9754);
and G8107 (W6710, W9755, W9756);
and G8108 (W6711, W9753, W9757);
and G8109 (W6712, W9758, W9759);
and G8110 (W6713, W9753, W9760);
and G8111 (W6714, W9761, W9762);
nor G8112 (W6715, W9763, W9764, W9765);
nor G8113 (W6716, W9766, W9767, W9768);
not G8114 (W6717, I320);
not G8115 (W6718, I321);
not G8116 (W6719, I322);
nor G8117 (W6720, W9769, W9770, W9771);
not G8118 (W6721, I323);
not G8119 (W6722, I324);
not G8120 (W6723, I325);
nor G8121 (W6724, W9772, W9773, W9774);
not G8122 (W6725, I326);
not G8123 (W6726, I327);
not G8124 (W6727, I328);
nor G8125 (W6728, W9775, W9776, W9777);
not G8126 (W6729, I329);
not G8127 (W6730, I330);
not G8128 (W6731, I331);
and G8129 (W6732, W9778, W9779);
and G8130 (W6733, W9780, W9781);
and G8131 (W6734, W9782, W9783);
and G8132 (W6735, W9784, W9785);
and G8133 (W6736, W9786, W9787);
and G8134 (W6737, W9788, W9789);
and G8135 (W6738, W9790, W9791);
and G8136 (W6739, W9792, W9793);
and G8137 (W6740, W9794, W9795);
and G8138 (W6741, W9796, W9797);
and G8139 (W6742, W9798, W9799);
and G8140 (W6743, W9800, W9801);
and G8141 (W6744, W9802, W9803);
and G8142 (W6745, W9804, W9805);
and G8143 (W6746, W9806, W9807);
and G8144 (W6747, W9808, W9809);
and G8145 (W6748, W9810, W9811);
and G8146 (W6749, W9812, W9813);
and G8147 (W6750, W9814, W9815);
and G8148 (W6751, W9816, W9817);
and G8149 (W6752, W9778, W9818);
and G8150 (W6753, W9819, W9820);
and G8151 (W6754, W9778, W9821);
and G8152 (W6755, W9822, W9823);
and G8153 (W6756, W9782, W9824);
and G8154 (W6757, W9825, W9826);
and G8155 (W6758, W9782, W9827);
and G8156 (W6759, W9828, W9829);
and G8157 (W6760, W9786, W9830);
and G8158 (W6761, W9831, W9832);
and G8159 (W6762, W9786, W9833);
and G8160 (W6763, W9834, W9835);
and G8161 (W6764, W9790, W9836);
and G8162 (W6765, W9837, W9838);
and G8163 (W6766, W9790, W9839);
and G8164 (W6767, W9840, W9841);
and G8165 (W6768, W9794, W9842);
and G8166 (W6769, W9843, W9844);
and G8167 (W6770, W9794, W9845);
and G8168 (W6771, W9846, W9847);
and G8169 (W6772, W9798, W9848);
and G8170 (W6773, W9849, W9850);
and G8171 (W6774, W9798, W9851);
and G8172 (W6775, W9852, W9853);
and G8173 (W6776, W9802, W9854);
and G8174 (W6777, W9855, W9856);
and G8175 (W6778, W9806, W9857);
and G8176 (W6779, W9858, W9859);
and G8177 (W6780, W9802, W9860);
and G8178 (W6781, W9861, W9862);
and G8179 (W6782, W9810, W9863);
and G8180 (W6783, W9864, W9865);
and G8181 (W6784, W9806, W9866);
and G8182 (W6785, W9867, W9868);
and G8183 (W6786, W9814, W9869);
and G8184 (W6787, W9870, W9871);
and G8185 (W6788, W9810, W9872);
and G8186 (W6789, W9873, W9874);
and G8187 (W6790, W9814, W9875);
and G8188 (W6791, W9876, W9877);
nor G8189 (W6792, W9878, W9879);
and G8190 (W6793, W9880, W9881, W9882);
nor G8191 (W6794, W9883, W9884);
nor G8192 (W6795, W9885, W9886);
nor G8193 (W6796, W9887, W9888);
nor G8194 (W6797, W9889, W9890);
nor G8195 (W6798, W9891, W9892);
nor G8196 (W6799, W9893, W9894);
nor G8197 (W6800, W9895, W9896);
nor G8198 (W6801, W9897, W9898);
nor G8199 (W6802, W9899, W9900);
not G8200 (W6803, I96);
and G8201 (W6804, W9901, W9902);
and G8202 (W6805, W9903, W9904);
and G8203 (W6806, W9901, W9905);
and G8204 (W6807, W9906, W9907);
and G8205 (W6808, W9901, W9908);
and G8206 (W6809, W9909, W9910);
and G8207 (W6810, W9806, W9911);
and G8208 (W6811, W9912, W9913);
and G8209 (W6812, W9806, W9914);
and G8210 (W6813, W9915, W9916);
and G8211 (W6814, W9806, W9917);
and G8212 (W6815, W9918, W9919);
and G8213 (W6816, W9814, W9920);
and G8214 (W6817, W9921, W9922);
and G8215 (W6818, W9814, W9923);
and G8216 (W6819, W9924, W9925);
and G8217 (W6820, W9814, W9926);
and G8218 (W6821, W9927, W9928);
and G8219 (W6822, W9929, W9930);
and G8220 (W6823, W9931, W9932);
and G8221 (W6824, W9929, W9933);
and G8222 (W6825, W9934, W9935);
and G8223 (W6826, W9929, W9936);
and G8224 (W6827, W9937, W9938);
nor G8225 (W6828, W9939, W9940);
nor G8226 (W6829, W9941, W9942);
nor G8227 (W6830, W9943, W9944);
nor G8228 (W6831, W9945, W9946);
nor G8229 (W6832, W9947, W9948);
nor G8230 (W6833, W9949, W9950, W9951);
nor G8231 (W6834, W9952, W9953);
nor G8232 (W6835, W9954, W9955);
nor G8233 (W6836, W9956, W9957);
and G8234 (W6837, W9958, W9959);
and G8235 (W6838, W9960, W9961);
and G8236 (W6839, W9958, W9962);
and G8237 (W6840, W9963, W9964);
and G8238 (W6841, W9958, W9965);
and G8239 (W6842, W9966, W9967);
and G8240 (W6843, W9968, W9969);
and G8241 (W6844, W9970, W9971);
and G8242 (W6845, W9968, W9972);
and G8243 (W6846, W9973, W9974);
and G8244 (W6847, W9968, W9975);
and G8245 (W6848, W9976, W9977);
and G8246 (W6849, W9978, W9979);
and G8247 (W6850, W9980, W9981);
and G8248 (W6851, W9978, W9982);
and G8249 (W6852, W9983, W9984);
and G8250 (W6853, W9978, W9985);
and G8251 (W6854, W9986, W9987);
and G8252 (W6855, W9988, W9989);
and G8253 (W6856, W9990, W9991);
and G8254 (W6857, W9988, W9992);
and G8255 (W6858, W9993, W9994);
and G8256 (W6859, W9988, W9995);
and G8257 (W6860, W9996, W9997);
and G8258 (W6861, I332, W9998);
and G8259 (W6862, W9999, W10000);
and G8260 (W6863, I332, W10001);
and G8261 (W6864, W10002, W10003);
and G8262 (W6865, I332, W10004);
and G8263 (W6866, W10005, W10006);
and G8264 (W6867, I333, W10007);
and G8265 (W6868, W10008, W10009);
and G8266 (W6869, I333, W10010);
and G8267 (W6870, W10011, W10012);
and G8268 (W6871, I333, W10013);
and G8269 (W6872, W10014, W10015);
and G8270 (W6873, I334, W10016);
and G8271 (W6874, W10017, W10018);
and G8272 (W6875, I334, W10019);
and G8273 (W6876, W10020, W10021);
and G8274 (W6877, I334, W10022);
and G8275 (W6878, W10023, W10024);
and G8276 (W6879, I335, W10025);
and G8277 (W6880, W10026, W10027);
and G8278 (W6881, I335, W10028);
and G8279 (W6882, W10029, W10030);
and G8280 (W6883, I335, W10031);
and G8281 (W6884, W10032, W10033);
and G8282 (W6885, I336, W10034);
and G8283 (W6886, W10035, W10036);
and G8284 (W6887, I336, W10037);
and G8285 (W6888, W10038, W10039);
and G8286 (W6889, I336, W10040);
and G8287 (W6890, W10041, W10042);
and G8288 (W6891, I337, W10043);
and G8289 (W6892, W10044, W10045);
and G8290 (W6893, I337, W10046);
and G8291 (W6894, W10047, W10048);
and G8292 (W6895, I337, W10049);
and G8293 (W6896, W10050, W10051);
and G8294 (W6897, I338, W10052);
and G8295 (W6898, W10053, W10054);
and G8296 (W6899, I338, W10055);
and G8297 (W6900, W10056, W10057);
and G8298 (W6901, I338, W10058);
and G8299 (W6902, W10059, W10060);
and G8300 (W6903, I339, W10061);
and G8301 (W6904, W10062, W10063);
and G8302 (W6905, I339, W10064);
and G8303 (W6906, W10065, W10066);
and G8304 (W6907, I339, W10067);
and G8305 (W6908, W10068, W10069);
and G8306 (W6909, I340, W10070);
and G8307 (W6910, W10071, W10072);
and G8308 (W6911, I340, W10073);
and G8309 (W6912, W10074, W10075);
and G8310 (W6913, I340, W10076);
and G8311 (W6914, W10077, W10078);
and G8312 (W6915, I341, W10079);
and G8313 (W6916, W10080, W10081);
and G8314 (W6917, I341, W10082);
and G8315 (W6918, W10083, W10084);
and G8316 (W6919, I341, W10085);
and G8317 (W6920, W10086, W10087);
nor G8318 (W6921, W10088, W10089);
and G8319 (W6922, W9958, W10090);
nor G8320 (W6923, W10091, W10092);
nor G8321 (W6924, W10093, W10094);
nor G8322 (W6925, W10095, W10096);
nor G8323 (W6926, W10097, W10098);
nor G8324 (W6927, W10099, W10100);
nor G8325 (W6928, W10101, W10102);
nor G8326 (W6929, W10103, W10104);
nor G8327 (W6930, W10105, W10106);
nor G8328 (W6931, W10107, W10108);
and G8329 (W6932, W10109, W10110);
and G8330 (W6933, W10111, W10112);
and G8331 (W6934, W10113, W10114);
and G8332 (W6935, W10115, W10116);
and G8333 (W6936, W10117, W10118);
and G8334 (W6937, W10119, W10120);
and G8335 (W6938, W10121, W10122);
and G8336 (W6939, W10123, W10124);
and G8337 (W6940, W10125, W10126);
and G8338 (W6941, W10127, W10128);
and G8339 (W6942, W10129, W10130);
and G8340 (W6943, W10131, W10132);
and G8341 (W6944, W10133, W10134);
and G8342 (W6945, W10135, W10136);
and G8343 (W6946, W10137, W10138);
and G8344 (W6947, W10135, W10139);
and G8345 (W6948, W10140, W10141);
and G8346 (W6949, W10135, W10142);
nor G8347 (W6950, W10143, W10144, W10145);
nor G8348 (W6951, W10146, W10147, W10148);
nor G8349 (W6952, W10149, W10150, W10151);
nor G8350 (W6953, W10152, W10153, W10154);
and G8351 (W6954, W10155, W10156);
and G8352 (W6955, W10157, W10158);
and G8353 (W6956, W10159, W10160);
and G8354 (W6957, W10157, W10161);
and G8355 (W6958, W10162, W10163);
and G8356 (W6959, W10157, W10164);
and G8357 (W6960, W10165, W10166);
and G8358 (W6961, W10167, W10168);
and G8359 (W6962, W10169, W10170);
and G8360 (W6963, W10167, W10171);
and G8361 (W6964, W10172, W10173);
and G8362 (W6965, W10167, W10174);
and G8363 (W6966, W10175, W10176);
and G8364 (W6967, W10177, W10178);
and G8365 (W6968, W10179, W10180);
and G8366 (W6969, W10181, W10182);
and G8367 (W6970, W10183, W10184);
and G8368 (W6971, W10181, W10185);
and G8369 (W6972, W10186, W10187);
and G8370 (W6973, W10181, W10188);
not G8371 (W6974, I342);
and G8372 (W6975, W10189, W10190);
and G8373 (W6976, W10191, W10192);
not G8374 (W6977, I343);
and G8375 (W6978, W10193, W10194);
and G8376 (W6979, W10191, W10195);
not G8377 (W6980, I344);
and G8378 (W6981, W10196, W10197);
and G8379 (W6982, W10191, W10198);
not G8380 (W6983, W10199);
and G8381 (W6984, W10200, W10201);
and G8382 (W6985, W10202, W10203);
and G8383 (W6986, W10204, W10205);
and G8384 (W6987, W10202, W10206);
and G8385 (W6988, W10207, W10208);
and G8386 (W6989, W10202, W10209);
not G8387 (W6990, W10210);
and G8388 (W6991, W10211, W10212);
and G8389 (W6992, W10213, W10214);
and G8390 (W6993, W10215, W10216);
and G8391 (W6994, W10213, W10217);
and G8392 (W6995, W10218, W10219);
and G8393 (W6996, W10213, W10220);
not G8394 (W6997, I345);
and G8395 (W6998, W10221, W10222);
and G8396 (W6999, W10223, W10224);
not G8397 (W7000, I346);
and G8398 (W7001, W10225, W10226);
and G8399 (W7002, W10223, W10227);
and G8400 (W7003, W10228, W10229);
and G8401 (W7004, W10223, W10230);
not G8402 (W7005, I347);
not G8403 (W7006, W10231);
and G8404 (W7007, W10232, W10233);
and G8405 (W7008, W10234, W10235);
and G8406 (W7009, W10236, W10237);
and G8407 (W7010, W10234, W10238);
and G8408 (W7011, W10239, W10240);
and G8409 (W7012, W10234, W10241);
and G8410 (W7013, W10242, I348);
and G8411 (W7014, W10243, I349);
and G8412 (W7015, W10244, I350);
and G8413 (W7016, W10242, I351);
and G8414 (W7017, W10243, I352);
and G8415 (W7018, W10244, I353);
and G8416 (W7019, W10245, W10246);
and G8417 (W7020, W10247, W10248);
and G8418 (W7021, W10247, W10249);
and G8419 (W7022, I354, W10250);
and G8420 (W7023, W10251, W10252);
and G8421 (W7024, I355, W10253);
and G8422 (W7025, W10254, W10255);
and G8423 (W7026, W10256, W10257);
and G8424 (W7027, W10258, W10259);
and G8425 (W7028, W10260, W10261);
and G8426 (W7029, W10262, W10263);
and G8427 (W7030, W10264, W10265);
and G8428 (W7031, W10266, W10267);
and G8429 (W7032, W10268, W10269);
and G8430 (W7033, W10270, W10271);
and G8431 (W7034, W10272, W10273);
not G8432 (W7035, W10274);
not G8433 (W7036, W10275);
not G8434 (W7037, W10276);
not G8435 (W7038, W10277);
not G8436 (W7039, W10278);
not G8437 (W7040, W10279);
not G8438 (W7041, W10280);
not G8439 (W7042, W10281);
not G8440 (W7043, W10282);
not G8441 (W7044, W10283);
and G8442 (W7045, W10284, W10285);
and G8443 (W7046, W10286, W10287);
and G8444 (W7047, W10284, W10288);
and G8445 (W7048, W10289, W10290);
and G8446 (W7049, W10284, W10291);
and G8447 (W7050, W10292, W10293);
and G8448 (W7051, W10294, W10295);
and G8449 (W7052, W10296, W10297);
and G8450 (W7053, W10298, W10299);
and G8451 (W7054, W10296, W10300);
and G8452 (W7055, W10301, W10302);
and G8453 (W7056, W10296, W10303);
and G8454 (W7057, W10304, W10305);
and G8455 (W7058, W10306, W10307);
and G8456 (W7059, W10308, W10309);
and G8457 (W7060, W10306, W10310);
and G8458 (W7061, W10311, W10312);
and G8459 (W7062, W10306, W10313);
and G8460 (W7063, W10314, W10315);
and G8461 (W7064, W10316, W10317);
and G8462 (W7065, W10318, W10319);
and G8463 (W7066, W10316, W10320);
and G8464 (W7067, W10321, W10322);
and G8465 (W7068, W10316, W10323);
and G8466 (W7069, W10324, W10325);
and G8467 (W7070, W10326, W10327);
and G8468 (W7071, W10328, W10329);
and G8469 (W7072, W10326, W10330);
and G8470 (W7073, W10331, W10332);
and G8471 (W7074, W10326, W10333);
and G8472 (W7075, W10334, W10335);
and G8473 (W7076, W10336, W10337);
and G8474 (W7077, W10338, W10339);
and G8475 (W7078, W10336, W10340);
and G8476 (W7079, W10341, W10342);
and G8477 (W7080, W10336, W10343);
and G8478 (W7081, W10344, W10345);
and G8479 (W7082, W10346, W10347);
and G8480 (W7083, W10348, W10349);
and G8481 (W7084, W10346, W10350);
and G8482 (W7085, W10351, W10352);
and G8483 (W7086, W10346, W10353);
and G8484 (W7087, W10354, W10355);
and G8485 (W7088, W10356, W10357);
and G8486 (W7089, W10358, W10359);
and G8487 (W7090, W10356, W10360);
and G8488 (W7091, W10361, W10362);
and G8489 (W7092, W10356, W10363);
and G8490 (W7093, W10364, W10365);
and G8491 (W7094, W10366, W10367);
and G8492 (W7095, W10368, W10369);
and G8493 (W7096, W10366, W10370);
and G8494 (W7097, W10371, W10372);
and G8495 (W7098, W10366, W10373);
and G8496 (W7099, W10374, W10375);
and G8497 (W7100, W10376, W10377);
and G8498 (W7101, W10378, W10379);
and G8499 (W7102, W10376, W10380);
and G8500 (W7103, W10381, W10382);
and G8501 (W7104, W10376, W10383);
and G8502 (W7105, W10384, W10385);
and G8503 (W7106, W10386, W10387);
and G8504 (W7107, W10388, W10389);
and G8505 (W7108, W10386, W10390);
and G8506 (W7109, W10391, W10392);
and G8507 (W7110, W10386, W10393);
and G8508 (W7111, W10394, W10395);
and G8509 (W7112, W10396, W10397);
and G8510 (W7113, W10398, W10399);
and G8511 (W7114, W10396, W10400);
and G8512 (W7115, W10401, W10402);
and G8513 (W7116, W10396, W10403);
and G8514 (W7117, W10404, W10405);
and G8515 (W7118, W10406, W10407);
and G8516 (W7119, W10408, W10409);
and G8517 (W7120, W10406, W10410);
and G8518 (W7121, W10411, W10412);
and G8519 (W7122, W10406, W10413);
and G8520 (W7123, W10414, W10415);
and G8521 (W7124, W10416, W10417);
and G8522 (W7125, W10418, W10419);
and G8523 (W7126, W10416, W10420);
and G8524 (W7127, W10421, W10422);
and G8525 (W7128, W10416, W10423);
and G8526 (W7129, W10424, W10425);
and G8527 (W7130, W10426, W10427);
and G8528 (W7131, W10424, W10428);
and G8529 (W7132, W10429, W10430);
and G8530 (W7133, W10424, W10431);
and G8531 (W7134, W10432, W10433);
not G8532 (W7135, W10434);
not G8533 (W7136, W10435);
and G8534 (W7137, W10436, W10437);
and G8535 (W7138, W10438, W10439);
and G8536 (W7139, W10440, W10441);
and G8537 (W7140, W10442, W10443);
and G8538 (W7141, W10444, W10445);
and G8539 (W7142, W10446, W10447);
and G8540 (W7143, W10448, W10449);
and G8541 (W7144, W10450, W10451);
and G8542 (W7145, W10436, W10452);
and G8543 (W7146, W10453, W10454);
and G8544 (W7147, W10436, W10455);
and G8545 (W7148, W10456, W10457);
and G8546 (W7149, W10440, W10458);
and G8547 (W7150, W10459, W10460);
and G8548 (W7151, W10440, W10461);
and G8549 (W7152, W10462, W10463);
and G8550 (W7153, W10444, W10464);
and G8551 (W7154, W10465, W10466);
and G8552 (W7155, W10444, W10467);
and G8553 (W7156, W10468, W10469);
and G8554 (W7157, W10448, W10470);
and G8555 (W7158, W10471, W10472);
and G8556 (W7159, W10448, W10473);
and G8557 (W7160, W10474, W10475);
and G8558 (W7161, W10476, W10477);
and G8559 (W7162, W10478, W10479);
and G8560 (W7163, W10480, W10481);
and G8561 (W7164, W10478, W10482);
and G8562 (W7165, W10483, W10484);
and G8563 (W7166, W10478, W10485);
and G8564 (W7167, W10486, W10487);
and G8565 (W7168, W10488, W10489);
and G8566 (W7169, W10486, W10490);
and G8567 (W7170, W10491, W10492);
and G8568 (W7171, W10486, W10493);
and G8569 (W7172, W10494, W10495);
and G8570 (W7173, W10496, W10497);
and G8571 (W7174, W10498, W10499);
and G8572 (W7175, W10500, W10501);
and G8573 (W7176, W10498, W10502);
and G8574 (W7177, W10503, W10504);
and G8575 (W7178, W10498, W10505);
and G8576 (W7179, W10506, W10507);
and G8577 (W7180, W10508, W10509);
and G8578 (W7181, W10510, W10511);
and G8579 (W7182, W10508, W10512);
and G8580 (W7183, W10513, W10514);
and G8581 (W7184, W10508, W10515);
and G8582 (W7185, W10516, W10517);
and G8583 (W7186, W10518, W10519);
and G8584 (W7187, W10520, W10521);
and G8585 (W7188, W10518, W10522);
and G8586 (W7189, W10523, W10524);
and G8587 (W7190, W10518, W10525);
and G8588 (W7191, W10526, W10527);
and G8589 (W7192, W10528, W10529);
and G8590 (W7193, W10526, W10530);
and G8591 (W7194, W10531, W10532);
and G8592 (W7195, W10526, W10533);
and G8593 (W7196, W10534, W10535);
nor G8594 (W7197, W10536, W10537, W10538);
nor G8595 (W7198, W10539, W10540, W10541);
not G8596 (W7199, I356);
not G8597 (W7200, I357);
not G8598 (W7201, I358);
nor G8599 (W7202, W10542, W10543, W10544);
not G8600 (W7203, I359);
not G8601 (W7204, I360);
not G8602 (W7205, I361);
nor G8603 (W7206, W10545, W10546, W10547);
not G8604 (W7207, I362);
not G8605 (W7208, I363);
not G8606 (W7209, I364);
nor G8607 (W7210, W10548, W10549, W10550);
not G8608 (W7211, I365);
not G8609 (W7212, I366);
not G8610 (W7213, I367);
and G8611 (W7214, W10551, W10552);
and G8612 (W7215, W10553, W10554);
and G8613 (W7216, W10555, W10556);
and G8614 (W7217, W10557, W10558);
and G8615 (W7218, W10559, W10560);
and G8616 (W7219, W10561, W10562);
and G8617 (W7220, W10563, W10564);
and G8618 (W7221, W10565, W10566);
and G8619 (W7222, W10567, W10568);
and G8620 (W7223, W10569, W10570);
and G8621 (W7224, W10571, W10572);
and G8622 (W7225, W10573, W10574);
and G8623 (W7226, W10575, W10576);
and G8624 (W7227, W10577, W10578);
and G8625 (W7228, W10579, W10580);
and G8626 (W7229, W10581, W10582);
and G8627 (W7230, W10583, W10584);
and G8628 (W7231, W10585, W10586);
and G8629 (W7232, W10587, W10588);
and G8630 (W7233, W10589, W10590);
and G8631 (W7234, W10587, W10591);
and G8632 (W7235, W10592, W10593);
and G8633 (W7236, W10551, W10594);
and G8634 (W7237, W10595, W10596);
and G8635 (W7238, W10551, W10597);
and G8636 (W7239, W10598, W10599);
and G8637 (W7240, W10555, W10600);
and G8638 (W7241, W10601, W10602);
and G8639 (W7242, W10555, W10603);
and G8640 (W7243, W10604, W10605);
and G8641 (W7244, W10559, W10606);
and G8642 (W7245, W10607, W10608);
and G8643 (W7246, W10559, W10609);
and G8644 (W7247, W10610, W10611);
and G8645 (W7248, W10563, W10612);
and G8646 (W7249, W10613, W10614);
and G8647 (W7250, W10563, W10615);
and G8648 (W7251, W10616, W10617);
and G8649 (W7252, W10567, W10618);
and G8650 (W7253, W10619, W10620);
and G8651 (W7254, W10567, W10621);
and G8652 (W7255, W10622, W10623);
and G8653 (W7256, W10571, W10624);
and G8654 (W7257, W10625, W10626);
and G8655 (W7258, W10575, W10627);
and G8656 (W7259, W10628, W10629);
and G8657 (W7260, W10571, W10630);
and G8658 (W7261, W10631, W10632);
and G8659 (W7262, W10579, W10633);
and G8660 (W7263, W10634, W10635);
and G8661 (W7264, W10575, W10636);
and G8662 (W7265, W10637, W10638);
and G8663 (W7266, W10583, W10639);
and G8664 (W7267, W10640, W10641);
and G8665 (W7268, W10579, W10642);
and G8666 (W7269, W10643, W10644);
and G8667 (W7270, W10583, W10645);
and G8668 (W7271, W10646, W10647);
and G8669 (W7272, W10587, W10648);
and G8670 (W7273, W10649, W10650);
nor G8671 (W7274, W10651, W10652);
and G8672 (W7275, W10653, W10654, W10655);
nor G8673 (W7276, W10656, W10657);
nor G8674 (W7277, W10658, W10659);
nor G8675 (W7278, W10660, W10661);
nor G8676 (W7279, W10662, W10663);
nor G8677 (W7280, W10664, W10665);
nor G8678 (W7281, W10666, W10667);
nor G8679 (W7282, W10668, W10669);
nor G8680 (W7283, W10670, W10671);
nor G8681 (W7284, W10672, W10673);
not G8682 (W7285, I145);
and G8683 (W7286, W10674, W10675);
and G8684 (W7287, W10676, W10677);
and G8685 (W7288, W10674, W10678);
and G8686 (W7289, W10679, W10680);
and G8687 (W7290, W10674, W10681);
and G8688 (W7291, W10682, W10683);
and G8689 (W7292, W10575, W10684);
and G8690 (W7293, W10685, W10686);
and G8691 (W7294, W10575, W10687);
and G8692 (W7295, W10688, W10689);
and G8693 (W7296, W10575, W10690);
and G8694 (W7297, W10691, W10692);
and G8695 (W7298, W10583, W10693);
and G8696 (W7299, W10694, W10695);
and G8697 (W7300, W10583, W10696);
and G8698 (W7301, W10697, W10698);
and G8699 (W7302, W10583, W10699);
and G8700 (W7303, W10700, W10701);
and G8701 (W7304, W10702, W10703);
and G8702 (W7305, W10704, W10705);
and G8703 (W7306, W10702, W10706);
and G8704 (W7307, W10707, W10708);
and G8705 (W7308, W10702, W10709);
and G8706 (W7309, W10710, W10711);
nor G8707 (W7310, W10712, W10713);
nor G8708 (W7311, W10714, W10715);
nor G8709 (W7312, W10716, W10717);
nor G8710 (W7313, W10718, W10719);
nor G8711 (W7314, W10720, W10721);
nor G8712 (W7315, W10722, W10723, W10724);
nor G8713 (W7316, W10725, W10726);
nor G8714 (W7317, W10727, W10728);
nor G8715 (W7318, W10729, W10730);
and G8716 (W7319, W10731, W10732);
and G8717 (W7320, W10733, W10734);
and G8718 (W7321, W10731, W10735);
and G8719 (W7322, W10736, W10737);
and G8720 (W7323, W10731, W10738);
and G8721 (W7324, W10739, W10740);
and G8722 (W7325, W10741, W10742);
and G8723 (W7326, W10743, W10744);
and G8724 (W7327, W10741, W10745);
and G8725 (W7328, W10746, W10747);
and G8726 (W7329, W10741, W10748);
and G8727 (W7330, W10749, W10750);
and G8728 (W7331, W10751, W10752);
and G8729 (W7332, W10753, W10754);
and G8730 (W7333, W10751, W10755);
and G8731 (W7334, W10756, W10757);
and G8732 (W7335, W10751, W10758);
and G8733 (W7336, W10759, W10760);
and G8734 (W7337, W10761, W10762);
and G8735 (W7338, W10763, W10764);
and G8736 (W7339, W10761, W10765);
and G8737 (W7340, W10766, W10767);
and G8738 (W7341, W10761, W10768);
and G8739 (W7342, W10769, W10770);
and G8740 (W7343, I368, W10771);
and G8741 (W7344, W10772, W10773);
and G8742 (W7345, I368, W10774);
and G8743 (W7346, W10775, W10776);
and G8744 (W7347, I368, W10777);
and G8745 (W7348, W10778, W10779);
and G8746 (W7349, I369, W10780);
and G8747 (W7350, W10781, W10782);
and G8748 (W7351, I369, W10783);
and G8749 (W7352, W10784, W10785);
and G8750 (W7353, I369, W10786);
and G8751 (W7354, W10787, W10788);
and G8752 (W7355, I370, W10789);
and G8753 (W7356, W10790, W10791);
and G8754 (W7357, I370, W10792);
and G8755 (W7358, W10793, W10794);
and G8756 (W7359, I370, W10795);
and G8757 (W7360, W10796, W10797);
and G8758 (W7361, I371, W10798);
and G8759 (W7362, W10799, W10800);
and G8760 (W7363, I371, W10801);
and G8761 (W7364, W10802, W10803);
and G8762 (W7365, I371, W10804);
and G8763 (W7366, W10805, W10806);
and G8764 (W7367, I372, W10807);
and G8765 (W7368, W10808, W10809);
and G8766 (W7369, I372, W10810);
and G8767 (W7370, W10811, W10812);
and G8768 (W7371, I372, W10813);
and G8769 (W7372, W10814, W10815);
and G8770 (W7373, I373, W10816);
and G8771 (W7374, W10817, W10818);
and G8772 (W7375, I373, W10819);
and G8773 (W7376, W10820, W10821);
and G8774 (W7377, I373, W10822);
and G8775 (W7378, W10823, W10824);
and G8776 (W7379, I374, W10825);
and G8777 (W7380, W10826, W10827);
and G8778 (W7381, I374, W10828);
and G8779 (W7382, W10829, W10830);
and G8780 (W7383, I374, W10831);
and G8781 (W7384, W10832, W10833);
and G8782 (W7385, I375, W10834);
and G8783 (W7386, W10835, W10836);
and G8784 (W7387, I375, W10837);
and G8785 (W7388, W10838, W10839);
and G8786 (W7389, I375, W10840);
and G8787 (W7390, W10841, W10842);
and G8788 (W7391, I376, W10843);
and G8789 (W7392, W10844, W10845);
and G8790 (W7393, I376, W10846);
and G8791 (W7394, W10847, W10848);
and G8792 (W7395, I376, W10849);
and G8793 (W7396, W10850, W10851);
and G8794 (W7397, I377, W10852);
and G8795 (W7398, W10853, W10854);
and G8796 (W7399, I377, W10855);
and G8797 (W7400, W10856, W10857);
and G8798 (W7401, I377, W10858);
and G8799 (W7402, W10859, W10860);
nor G8800 (W7403, W10861, W10862);
and G8801 (W7404, W10731, W10863);
nor G8802 (W7405, W10864, W10865);
nor G8803 (W7406, W10866, W10867);
nor G8804 (W7407, W10868, W10869);
nor G8805 (W7408, W10870, W10871);
nor G8806 (W7409, W10872, W10873);
nor G8807 (W7410, W10874, W10875);
nor G8808 (W7411, W10876, W10877);
nor G8809 (W7412, W10878, W10879);
nor G8810 (W7413, W10880, W10881);
and G8811 (W7414, W10882, W10883);
and G8812 (W7415, W10884, W10885);
and G8813 (W7416, W10886, W10887);
and G8814 (W7417, W10888, W10889);
and G8815 (W7418, W10890, W10891);
and G8816 (W7419, W10892, W10893);
and G8817 (W7420, W10894, W10895);
and G8818 (W7421, W10896, W10897);
and G8819 (W7422, W10898, W10899);
and G8820 (W7423, W10900, W10901);
and G8821 (W7424, W10902, W10903);
and G8822 (W7425, W10904, W10905);
and G8823 (W7426, W10906, W10907);
and G8824 (W7427, W10908, W10909);
and G8825 (W7428, W10910, W10911);
and G8826 (W7429, W10908, W10912);
and G8827 (W7430, W10913, W10914);
and G8828 (W7431, W10908, W10915);
nor G8829 (W7432, W10916, W10917, W10918);
nor G8830 (W7433, W10919, W10920, W10921);
nor G8831 (W7434, W10922, W10923, W10924);
nor G8832 (W7435, W10925, W10926, W10927);
and G8833 (W7436, W10928, W10929);
and G8834 (W7437, W10930, W10931);
and G8835 (W7438, W10932, W10933);
and G8836 (W7439, W10930, W10934);
and G8837 (W7440, W10935, W10936);
and G8838 (W7441, W10930, W10937);
and G8839 (W7442, W10938, W10939);
and G8840 (W7443, W10940, W10941);
and G8841 (W7444, W10942, W10943);
and G8842 (W7445, W10940, W10944);
and G8843 (W7446, W10945, W10946);
and G8844 (W7447, W10940, W10947);
and G8845 (W7448, W10948, W10949);
and G8846 (W7449, W10950, W10951);
and G8847 (W7450, W10952, W10953);
and G8848 (W7451, W10954, W10955);
and G8849 (W7452, W10956, W10957);
and G8850 (W7453, W10954, W10958);
and G8851 (W7454, W10959, W10960);
and G8852 (W7455, W10954, W10961);
not G8853 (W7456, I378);
and G8854 (W7457, W10962, W10963);
and G8855 (W7458, W10964, W10965);
not G8856 (W7459, I379);
and G8857 (W7460, W10966, W10967);
and G8858 (W7461, W10964, W10968);
not G8859 (W7462, I380);
and G8860 (W7463, W10969, W10970);
and G8861 (W7464, W10964, W10971);
not G8862 (W7465, W10972);
and G8863 (W7466, W10973, W10974);
and G8864 (W7467, W10975, W10976);
and G8865 (W7468, W10977, W10978);
and G8866 (W7469, W10975, W10979);
and G8867 (W7470, W10980, W10981);
and G8868 (W7471, W10975, W10982);
not G8869 (W7472, W10983);
and G8870 (W7473, W10984, W10985);
and G8871 (W7474, W10986, W10987);
and G8872 (W7475, W10988, W10989);
and G8873 (W7476, W10986, W10990);
and G8874 (W7477, W10991, W10992);
and G8875 (W7478, W10986, W10993);
not G8876 (W7479, I381);
and G8877 (W7480, W10994, W10995);
and G8878 (W7481, W10996, W10997);
not G8879 (W7482, I382);
and G8880 (W7483, W10998, W10999);
and G8881 (W7484, W10996, W11000);
and G8882 (W7485, W11001, W11002);
and G8883 (W7486, W10996, W11003);
not G8884 (W7487, I383);
not G8885 (W7488, W11004);
and G8886 (W7489, W11005, W11006);
and G8887 (W7490, W11007, W11008);
and G8888 (W7491, W11009, W11010);
and G8889 (W7492, W11007, W11011);
and G8890 (W7493, W11012, W11013);
and G8891 (W7494, W11007, W11014);
and G8892 (W7495, W11015, I384);
and G8893 (W7496, W11016, I385);
and G8894 (W7497, W11017, I386);
and G8895 (W7498, W11015, I387);
and G8896 (W7499, W11016, I388);
and G8897 (W7500, W11017, I389);
and G8898 (W7501, W11018, W11019);
and G8899 (W7502, W11020, W11021);
and G8900 (W7503, W11020, W11022);
and G8901 (W7504, I390, W11023);
and G8902 (W7505, W11024, W11025);
and G8903 (W7506, I391, W11026);
and G8904 (W7507, W11027, W11028);
and G8905 (W7508, W11029, W11030);
and G8906 (W7509, W11031, W11032);
and G8907 (W7510, W11033, W11034);
and G8908 (W7511, W11035, W11036);
and G8909 (W7512, W11037, W11038);
and G8910 (W7513, W11039, W11040);
and G8911 (W7514, W11041, W11042);
and G8912 (W7515, W11043, W11044);
and G8913 (W7516, W11045, W11046);
not G8914 (W7517, W11047);
not G8915 (W7518, W11048);
not G8916 (W7519, W11049);
not G8917 (W7520, W11050);
not G8918 (W7521, W11051);
not G8919 (W7522, W11052);
not G8920 (W7523, W11053);
not G8921 (W7524, W11054);
not G8922 (W7525, W11055);
not G8923 (W7526, W11056);
and G8924 (W7527, W11057, W11058);
and G8925 (W7528, W11059, W11060);
and G8926 (W7529, W11057, W11061);
and G8927 (W7530, W11062, W11063);
and G8928 (W7531, W11057, W11064);
and G8929 (W7532, W11065, W11066);
and G8930 (W7533, W11067, W11068);
and G8931 (W7534, W11069, W11070);
and G8932 (W7535, W11071, W11072);
and G8933 (W7536, W11069, W11073);
and G8934 (W7537, W11074, W11075);
and G8935 (W7538, W11069, W11076);
and G8936 (W7539, W11077, W11078);
and G8937 (W7540, W11079, W11080);
and G8938 (W7541, W11081, W11082);
and G8939 (W7542, W11079, W11083);
and G8940 (W7543, W11084, W11085);
and G8941 (W7544, W11079, W11086);
and G8942 (W7545, W11087, W11088);
and G8943 (W7546, W11089, W11090);
and G8944 (W7547, W11091, W11092);
and G8945 (W7548, W11089, W11093);
and G8946 (W7549, W11094, W11095);
and G8947 (W7550, W11089, W11096);
and G8948 (W7551, W11097, W11098);
and G8949 (W7552, W11099, W11100);
and G8950 (W7553, W11101, W11102);
and G8951 (W7554, W11099, W11103);
and G8952 (W7555, W11104, W11105);
and G8953 (W7556, W11099, W11106);
and G8954 (W7557, W11107, W11108);
and G8955 (W7558, W11109, W11110);
and G8956 (W7559, W11111, W11112);
and G8957 (W7560, W11109, W11113);
and G8958 (W7561, W11114, W11115);
and G8959 (W7562, W11109, W11116);
and G8960 (W7563, W11117, W11118);
and G8961 (W7564, W11119, W11120);
and G8962 (W7565, W11121, W11122);
and G8963 (W7566, W11119, W11123);
and G8964 (W7567, W11124, W11125);
and G8965 (W7568, W11119, W11126);
and G8966 (W7569, W11127, W11128);
and G8967 (W7570, W11129, W11130);
and G8968 (W7571, W11131, W11132);
and G8969 (W7572, W11129, W11133);
and G8970 (W7573, W11134, W11135);
and G8971 (W7574, W11129, W11136);
and G8972 (W7575, W11137, W11138);
and G8973 (W7576, W11139, W11140);
and G8974 (W7577, W11141, W11142);
and G8975 (W7578, W11139, W11143);
and G8976 (W7579, W11144, W11145);
and G8977 (W7580, W11139, W11146);
and G8978 (W7581, W11147, W11148);
and G8979 (W7582, W11149, W11150);
and G8980 (W7583, W11151, W11152);
and G8981 (W7584, W11149, W11153);
and G8982 (W7585, W11154, W11155);
and G8983 (W7586, W11149, W11156);
and G8984 (W7587, W11157, W11158);
and G8985 (W7588, W11159, W11160);
and G8986 (W7589, W11161, W11162);
and G8987 (W7590, W11159, W11163);
and G8988 (W7591, W11164, W11165);
and G8989 (W7592, W11159, W11166);
and G8990 (W7593, W11167, W11168);
and G8991 (W7594, W11169, W11170);
and G8992 (W7595, W11171, W11172);
and G8993 (W7596, W11169, W11173);
and G8994 (W7597, W11174, W11175);
and G8995 (W7598, W11169, W11176);
and G8996 (W7599, W11177, W11178);
and G8997 (W7600, W11179, W11180);
and G8998 (W7601, W11181, W11182);
and G8999 (W7602, W11179, W11183);
and G9000 (W7603, W11184, W11185);
and G9001 (W7604, W11179, W11186);
and G9002 (W7605, W11187, W11188);
and G9003 (W7606, W11189, W11190);
and G9004 (W7607, W11191, W11192);
and G9005 (W7608, W11189, W11193);
and G9006 (W7609, W11194, W11195);
and G9007 (W7610, W11189, W11196);
and G9008 (W7611, W11197, W11198);
and G9009 (W7612, W11199, W11200);
and G9010 (W7613, W11197, W11201);
and G9011 (W7614, W11202, W11203);
and G9012 (W7615, W11197, W11204);
and G9013 (W7616, W11205, W11206);
not G9014 (W7617, W11207);
not G9015 (W7618, W11208);
and G9016 (W7619, W11209, W11210);
and G9017 (W7620, W11211, W11212);
and G9018 (W7621, W11213, W11214);
and G9019 (W7622, W11215, W11216);
and G9020 (W7623, W11217, W11218);
and G9021 (W7624, W11219, W11220);
and G9022 (W7625, W11221, W11222);
and G9023 (W7626, W11223, W11224);
and G9024 (W7627, W11209, W11225);
and G9025 (W7628, W11226, W11227);
and G9026 (W7629, W11209, W11228);
and G9027 (W7630, W11229, W11230);
and G9028 (W7631, W11213, W11231);
and G9029 (W7632, W11232, W11233);
and G9030 (W7633, W11213, W11234);
and G9031 (W7634, W11235, W11236);
and G9032 (W7635, W11217, W11237);
and G9033 (W7636, W11238, W11239);
and G9034 (W7637, W11217, W11240);
and G9035 (W7638, W11241, W11242);
and G9036 (W7639, W11221, W11243);
and G9037 (W7640, W11244, W11245);
and G9038 (W7641, W11221, W11246);
and G9039 (W7642, W11247, W11248);
and G9040 (W7643, W11249, W11250);
and G9041 (W7644, W11251, W11252);
and G9042 (W7645, W11253, W11254);
and G9043 (W7646, W11251, W11255);
and G9044 (W7647, W11256, W11257);
and G9045 (W7648, W11251, W11258);
and G9046 (W7649, W11259, W11260);
and G9047 (W7650, W11261, W11262);
and G9048 (W7651, W11259, W11263);
and G9049 (W7652, W11264, W11265);
and G9050 (W7653, W11259, W11266);
and G9051 (W7654, W11267, W11268);
and G9052 (W7655, W11269, W11270);
and G9053 (W7656, W11271, W11272);
and G9054 (W7657, W11273, W11274);
and G9055 (W7658, W11271, W11275);
and G9056 (W7659, W11276, W11277);
and G9057 (W7660, W11271, W11278);
and G9058 (W7661, W11279, W11280);
and G9059 (W7662, W11281, W11282);
and G9060 (W7663, W11283, W11284);
and G9061 (W7664, W11281, W11285);
and G9062 (W7665, W11286, W11287);
and G9063 (W7666, W11281, W11288);
and G9064 (W7667, W11289, W11290);
and G9065 (W7668, W11291, W11292);
and G9066 (W7669, W11293, W11294);
and G9067 (W7670, W11291, W11295);
and G9068 (W7671, W11296, W11297);
and G9069 (W7672, W11291, W11298);
and G9070 (W7673, W11299, W11300);
and G9071 (W7674, W11301, W11302);
and G9072 (W7675, W11299, W11303);
and G9073 (W7676, W11304, W11305);
and G9074 (W7677, W11299, W11306);
and G9075 (W7678, W11307, W11308);
nor G9076 (W7679, W11309, W11310, W11311);
nor G9077 (W7680, W11312, W11313, W11314);
not G9078 (W7681, I392);
not G9079 (W7682, I393);
not G9080 (W7683, I394);
nor G9081 (W7684, W11315, W11316, W11317);
not G9082 (W7685, I395);
not G9083 (W7686, I396);
not G9084 (W7687, I397);
nor G9085 (W7688, W11318, W11319, W11320);
not G9086 (W7689, I398);
not G9087 (W7690, I399);
not G9088 (W7691, I400);
nor G9089 (W7692, W11321, W11322, W11323);
not G9090 (W7693, I401);
not G9091 (W7694, I402);
not G9092 (W7695, I403);
and G9093 (W7696, W11324, W11325);
and G9094 (W7697, W11326, W11327);
and G9095 (W7698, W11328, W11329);
and G9096 (W7699, W11330, W11331);
and G9097 (W7700, W11332, W11333);
and G9098 (W7701, W11334, W11335);
and G9099 (W7702, W11336, W11337);
and G9100 (W7703, W11338, W11339);
and G9101 (W7704, W11340, W11341);
and G9102 (W7705, W11342, W11343);
and G9103 (W7706, W11344, W11345);
and G9104 (W7707, W11346, W11347);
and G9105 (W7708, W11348, W11349);
and G9106 (W7709, W11350, W11351);
and G9107 (W7710, W11352, W11353);
and G9108 (W7711, W11354, W11355);
and G9109 (W7712, W11356, W11357);
and G9110 (W7713, W11358, W11359);
and G9111 (W7714, W11356, W11360);
and G9112 (W7715, W11361, W11362);
and G9113 (W7716, W11363, W11364);
and G9114 (W7717, W11365, W11366);
and G9115 (W7718, W11363, W11367);
and G9116 (W7719, W11368, W11369);
and G9117 (W7720, W11324, W11370);
and G9118 (W7721, W11371, W11372);
and G9119 (W7722, W11324, W11373);
and G9120 (W7723, W11374, W11375);
and G9121 (W7724, W11328, W11376);
and G9122 (W7725, W11377, W11378);
and G9123 (W7726, W11328, W11379);
and G9124 (W7727, W11380, W11381);
and G9125 (W7728, W11332, W11382);
and G9126 (W7729, W11383, W11384);
and G9127 (W7730, W11332, W11385);
and G9128 (W7731, W11386, W11387);
and G9129 (W7732, W11336, W11388);
and G9130 (W7733, W11389, W11390);
and G9131 (W7734, W11336, W11391);
and G9132 (W7735, W11392, W11393);
and G9133 (W7736, W11340, W11394);
and G9134 (W7737, W11395, W11396);
and G9135 (W7738, W11344, W11397);
and G9136 (W7739, W11398, W11399);
and G9137 (W7740, W11340, W11400);
and G9138 (W7741, W11401, W11402);
and G9139 (W7742, W11348, W11403);
and G9140 (W7743, W11404, W11405);
and G9141 (W7744, W11344, W11406);
and G9142 (W7745, W11407, W11408);
and G9143 (W7746, W11352, W11409);
and G9144 (W7747, W11410, W11411);
and G9145 (W7748, W11348, W11412);
and G9146 (W7749, W11413, W11414);
and G9147 (W7750, W11352, W11415);
and G9148 (W7751, W11416, W11417);
and G9149 (W7752, W11356, W11418);
and G9150 (W7753, W11419, W11420);
and G9151 (W7754, W11363, W11421);
and G9152 (W7755, W11422, W11423);
nor G9153 (W7756, W11424, W11425);
and G9154 (W7757, W11426, W11427, W11428);
nor G9155 (W7758, W11429, W11430);
nor G9156 (W7759, W11431, W11432);
nor G9157 (W7760, W11433, W11434);
nor G9158 (W7761, W11435, W11436);
nor G9159 (W7762, W11437, W11438);
nor G9160 (W7763, W11439, W11440);
nor G9161 (W7764, W11441, W11442);
nor G9162 (W7765, W11443, W11444);
nor G9163 (W7766, W11445, W11446);
not G9164 (W7767, I194);
and G9165 (W7768, W11447, W11448);
and G9166 (W7769, W11449, W11450);
and G9167 (W7770, W11447, W11451);
and G9168 (W7771, W11452, W11453);
and G9169 (W7772, W11447, W11454);
and G9170 (W7773, W11455, W11456);
and G9171 (W7774, W11344, W11457);
and G9172 (W7775, W11458, W11459);
and G9173 (W7776, W11344, W11460);
and G9174 (W7777, W11461, W11462);
and G9175 (W7778, W11344, W11463);
and G9176 (W7779, W11464, W11465);
and G9177 (W7780, W11352, W11466);
and G9178 (W7781, W11467, W11468);
and G9179 (W7782, W11352, W11469);
and G9180 (W7783, W11470, W11471);
and G9181 (W7784, W11352, W11472);
and G9182 (W7785, W11473, W11474);
and G9183 (W7786, W11475, W11476);
and G9184 (W7787, W11477, W11478);
and G9185 (W7788, W11475, W11479);
and G9186 (W7789, W11480, W11481);
and G9187 (W7790, W11475, W11482);
and G9188 (W7791, W11483, W11484);
not G9189 (W7792, W11485);
not G9190 (W7793, W11486);
and G9191 (W7794, W11487, W11488);
and G9192 (W7795, W11489, W11490);
and G9193 (W7796, W7806, W11491);
and G9194 (W7797, W11489, W11492);
and G9195 (W7798, W7857, W11493);
and G9196 (W7799, W11494, W11495);
and G9197 (W7800, W11496, W11497);
and G9198 (W7801, W11494, W11498);
not G9199 (W7802, W11499);
not G9200 (W7803, W11500);
not G9201 (W7804, W11501);
not G9202 (W7805, W11502);
not G9203 (W7806, I404);
and G9204 (W7807, W11503, W11504);
and G9205 (W7808, W11505, W11506);
and G9206 (W7809, W11507, W11508);
and G9207 (W7810, W11509, W11510);
and G9208 (W7811, W11511, W11512);
and G9209 (W7812, W11513, W11514);
and G9210 (W7813, W11515, W11516);
and G9211 (W7814, W11517, W11518);
and G9212 (W7815, W11519, W11520);
and G9213 (W7816, W11521, W11522);
and G9214 (W7817, W11523, W11524);
and G9215 (W7818, W11525, W11526);
and G9216 (W7819, W11527, W11528);
and G9217 (W7820, W11529, W11530);
and G9218 (W7821, W11531, W11532);
and G9219 (W7822, W11533, W11534);
not G9220 (W7823, I405);
and G9221 (W7824, W11535, W11536);
and G9222 (W7825, W11537, W11538);
and G9223 (W7826, W11539, W11540);
and G9224 (W7827, W11541, W11542);
and G9225 (W7828, W11543, W11544);
and G9226 (W7829, W11545, W11546);
and G9227 (W7830, W11547, W11548);
and G9228 (W7831, W11549, W11550);
and G9229 (W7832, W11551, W11552);
and G9230 (W7833, W11553, W11554);
and G9231 (W7834, W11555, W11556);
and G9232 (W7835, W11557, W11558);
and G9233 (W7836, W11559, W11560);
and G9234 (W7837, W11561, W11562);
and G9235 (W7838, W11563, W11564);
and G9236 (W7839, W11565, W11566);
not G9237 (W7840, I406);
and G9238 (W7841, W11567, W11568);
and G9239 (W7842, W11505, W11569);
and G9240 (W7843, W11570, W11571);
and G9241 (W7844, W11509, W11572);
and G9242 (W7845, W11573, W11574);
and G9243 (W7846, W11513, W11575);
and G9244 (W7847, W11576, W11577);
and G9245 (W7848, W11517, W11578);
and G9246 (W7849, W11579, W11580);
and G9247 (W7850, W11521, W11581);
and G9248 (W7851, W11582, W11583);
and G9249 (W7852, W11525, W11584);
and G9250 (W7853, W11585, W11586);
and G9251 (W7854, W11529, W11587);
and G9252 (W7855, W11588, W11589);
and G9253 (W7856, W11533, W11590);
not G9254 (W7857, I407);
and G9255 (W7858, W11591, W11592);
and G9256 (W7859, W11537, W11593);
and G9257 (W7860, W11594, W11595);
and G9258 (W7861, W11541, W11596);
and G9259 (W7862, W11597, W11598);
and G9260 (W7863, W11545, W11599);
and G9261 (W7864, W11600, W11601);
and G9262 (W7865, W11549, W11602);
and G9263 (W7866, W11603, W11604);
and G9264 (W7867, W11553, W11605);
and G9265 (W7868, W11606, W11607);
and G9266 (W7869, W11557, W11608);
and G9267 (W7870, W11609, W11610);
and G9268 (W7871, W11561, W11611);
and G9269 (W7872, W11612, W11613);
and G9270 (W7873, W11565, W11614);
nand G9271 (W7874, I408, W11615);
nand G9272 (W7875, W11616, W11615);
nand G9273 (W7876, I409, W11617);
nand G9274 (W7877, W11618, W11617);
or G9275 (W7878, I410, W11619);
not G9276 (W7879, W11620);
not G9277 (W7880, W11620);
not G9278 (W7881, W11620);
not G9279 (W7882, W11620);
nor G9280 (W7883, W11621, W11622);
not G9281 (W7884, W7888);
nor G9282 (W7885, W11623, W11624);
nor G9283 (W7886, W11625, W11626);
nor G9284 (W7887, W11627, W11628);
nor G9285 (W7888, W11629, I411);
nor G9286 (W7889, W11630, W11631);
not G9287 (W7890, W7897);
nor G9288 (W7891, W11632, W11633);
nor G9289 (W7892, W11634, W11635);
nor G9290 (W7893, W11636, W11637);
nor G9291 (W7894, W11638, W11639);
nor G9292 (W7895, W11640, W11641);
nor G9293 (W7896, W11642, W11643);
nor G9294 (W7897, I411, W11644);
not G9295 (W7898, W11645);
not G9296 (W7899, I412);
not G9297 (W7900, W11646);
not G9298 (W7901, W11646);
not G9299 (W7902, W11646);
not G9300 (W7903, W11646);
not G9301 (W7904, W11646);
not G9302 (W7905, W11646);
not G9303 (W7906, W11646);
not G9304 (W7907, W11646);
not G9305 (W7908, W11646);
not G9306 (W7909, W11646);
not G9307 (W7910, W11646);
not G9308 (W7911, W11646);
not G9309 (W7912, I413);
not G9310 (W7913, W7898);
not G9311 (W7914, I414);
not G9312 (W7915, W11647);
not G9313 (W7916, W11648);
nand G9314 (W7917, W11649, W11650);
nand G9315 (W7918, W7919, W11650);
nand G9316 (W7919, W11651, W11652);
nand G9317 (W7920, W7919, W7921);
nor G9318 (W7921, W11653, W11654);
nand G9319 (W7922, W11655, W11656);
nand G9320 (W7923, W7924, W11656);
nand G9321 (W7924, W11657, W11658);
nand G9322 (W7925, W7924, W7921);
not G9323 (W7926, I415);
not G9324 (W7927, W7929);
not G9325 (W7928, I416);
not G9326 (W7929, W11659);
not G9327 (W7930, I417);
not G9328 (W7931, W7933);
not G9329 (W7932, I418);
not G9330 (W7933, W11660);
not G9331 (W7934, I419);
not G9332 (W7935, W7937);
not G9333 (W7936, I420);
not G9334 (W7937, W11661);
not G9335 (W7938, I421);
not G9336 (W7939, W7941);
not G9337 (W7940, I422);
not G9338 (W7941, W11662);
not G9339 (W7942, I423);
not G9340 (W7943, W7945);
not G9341 (W7944, I424);
not G9342 (W7945, W11663);
not G9343 (W7946, I425);
not G9344 (W7947, W7949);
not G9345 (W7948, I426);
not G9346 (W7949, W11664);
not G9347 (W7950, I427);
not G9348 (W7951, W7953);
not G9349 (W7952, I428);
not G9350 (W7953, W11665);
not G9351 (W7954, I429);
not G9352 (W7955, W7957);
not G9353 (W7956, I430);
not G9354 (W7957, W11666);
not G9355 (W7958, I431);
not G9356 (W7959, W7961);
not G9357 (W7960, I432);
not G9358 (W7961, W11667);
not G9359 (W7962, I433);
not G9360 (W7963, W7965);
not G9361 (W7964, I434);
not G9362 (W7965, W11668);
not G9363 (W7966, I435);
not G9364 (W7967, W7969);
not G9365 (W7968, I436);
not G9366 (W7969, W11669);
not G9367 (W7970, I437);
not G9368 (W7971, W7973);
not G9369 (W7972, I438);
not G9370 (W7973, W11670);
not G9371 (W7974, I439);
not G9372 (W7975, W7977);
not G9373 (W7976, I440);
not G9374 (W7977, W11671);
not G9375 (W7978, I441);
not G9376 (W7979, W7981);
not G9377 (W7980, I442);
not G9378 (W7981, W11672);
not G9379 (W7982, I443);
not G9380 (W7983, W7985);
not G9381 (W7984, I444);
not G9382 (W7985, W11673);
not G9383 (W7986, I445);
not G9384 (W7987, W7989);
not G9385 (W7988, I446);
not G9386 (W7989, W11674);
not G9387 (W7990, I447);
not G9388 (W7991, W7993);
not G9389 (W7992, I448);
not G9390 (W7993, W11675);
not G9391 (W7994, I449);
not G9392 (W7995, W7997);
not G9393 (W7996, I450);
not G9394 (W7997, W11676);
not G9395 (W7998, I451);
not G9396 (W7999, I1);
not G9397 (W8000, I390);
not G9398 (W8001, W8003);
not G9399 (W8002, W11677);
not G9400 (W8003, W11678);
not G9401 (W8004, I354);
not G9402 (W8005, W8007);
not G9403 (W8006, W11679);
not G9404 (W8007, W11680);
not G9405 (W8008, I318);
not G9406 (W8009, W8011);
not G9407 (W8010, W11681);
not G9408 (W8011, W11682);
not G9409 (W8012, I282);
not G9410 (W8013, W8015);
not G9411 (W8014, W11683);
not G9412 (W8015, W11684);
not G9413 (W8016, I452);
not G9414 (W8017, W8019);
not G9415 (W8018, W11685);
not G9416 (W8019, W11686);
not G9417 (W8020, I453);
not G9418 (W8021, W8022);
not G9419 (W8022, W11687);
not G9420 (W8023, I454);
not G9421 (W8024, W8025);
not G9422 (W8025, W11688);
not G9423 (W8026, I455);
not G9424 (W8027, W8029);
not G9425 (W8028, W11689);
not G9426 (W8029, W11690);
not G9427 (W8030, I456);
not G9428 (W8031, W8032);
not G9429 (W8032, W11691);
not G9430 (W8033, I457);
not G9431 (W8034, W8035);
not G9432 (W8035, W11692);
not G9433 (W8036, I458);
not G9434 (W8037, W8039);
not G9435 (W8038, W11693);
not G9436 (W8039, W11694);
not G9437 (W8040, I459);
not G9438 (W8041, W8042);
not G9439 (W8042, W11695);
not G9440 (W8043, I460);
not G9441 (W8044, W8045);
not G9442 (W8045, W11696);
not G9443 (W8046, I461);
not G9444 (W8047, W8049);
not G9445 (W8048, W11697);
not G9446 (W8049, W11698);
not G9447 (W8050, I462);
not G9448 (W8051, W8052);
not G9449 (W8052, W11699);
not G9450 (W8053, I463);
not G9451 (W8054, W8055);
not G9452 (W8055, W11700);
not G9453 (W8056, I464);
not G9454 (W8057, W8059);
not G9455 (W8058, W11701);
not G9456 (W8059, W11702);
not G9457 (W8060, I465);
not G9458 (W8061, W8062);
not G9459 (W8062, W11703);
not G9460 (W8063, I466);
not G9461 (W8064, W8065);
not G9462 (W8065, W11704);
not G9463 (W8066, I467);
not G9464 (W8067, W8069);
not G9465 (W8068, W11705);
not G9466 (W8069, W11706);
not G9467 (W8070, I468);
not G9468 (W8071, W8072);
not G9469 (W8072, W11707);
not G9470 (W8073, I469);
not G9471 (W8074, W8075);
not G9472 (W8075, W11708);
not G9473 (W8076, I470);
not G9474 (W8077, W8079);
not G9475 (W8078, W11709);
not G9476 (W8079, W11710);
not G9477 (W8080, I471);
not G9478 (W8081, W8082);
not G9479 (W8082, W11711);
not G9480 (W8083, I472);
not G9481 (W8084, W8085);
not G9482 (W8085, W11712);
not G9483 (W8086, I473);
not G9484 (W8087, W8089);
not G9485 (W8088, W11713);
not G9486 (W8089, W11714);
not G9487 (W8090, I474);
not G9488 (W8091, W8092);
not G9489 (W8092, W11715);
not G9490 (W8093, I475);
not G9491 (W8094, W8095);
not G9492 (W8095, W11716);
not G9493 (W8096, I476);
not G9494 (W8097, W8099);
not G9495 (W8098, W11717);
not G9496 (W8099, W11718);
not G9497 (W8100, I477);
not G9498 (W8101, W8102);
not G9499 (W8102, W11719);
not G9500 (W8103, I478);
not G9501 (W8104, W8105);
not G9502 (W8105, W11720);
not G9503 (W8106, I479);
not G9504 (W8107, W8109);
not G9505 (W8108, W11721);
not G9506 (W8109, W11722);
not G9507 (W8110, I480);
not G9508 (W8111, W8112);
not G9509 (W8112, W11723);
not G9510 (W8113, I481);
not G9511 (W8114, W8115);
not G9512 (W8115, W11724);
not G9513 (W8116, I482);
not G9514 (W8117, W8119);
not G9515 (W8118, W11725);
not G9516 (W8119, W11726);
not G9517 (W8120, I483);
not G9518 (W8121, W8122);
not G9519 (W8122, W11727);
not G9520 (W8123, I484);
not G9521 (W8124, W8125);
not G9522 (W8125, W11728);
not G9523 (W8126, I485);
not G9524 (W8127, W8129);
not G9525 (W8128, W11729);
not G9526 (W8129, W11730);
not G9527 (W8130, I486);
not G9528 (W8131, W8132);
not G9529 (W8132, W11731);
not G9530 (W8133, I487);
not G9531 (W8134, W8135);
not G9532 (W8135, W11732);
not G9533 (W8136, I488);
not G9534 (W8137, W8139);
not G9535 (W8138, W11733);
not G9536 (W8139, W11734);
not G9537 (W8140, I489);
not G9538 (W8141, W8142);
not G9539 (W8142, W11735);
not G9540 (W8143, I490);
not G9541 (W8144, W8145);
not G9542 (W8145, W11736);
not G9543 (W8146, I491);
not G9544 (W8147, W8149);
not G9545 (W8148, W11737);
not G9546 (W8149, W11738);
not G9547 (W8150, I492);
not G9548 (W8151, W8152);
not G9549 (W8152, W11739);
not G9550 (W8153, I493);
not G9551 (W8154, W8155);
not G9552 (W8155, W11740);
not G9553 (W8156, I494);
not G9554 (W8157, W8159);
not G9555 (W8158, W11741);
not G9556 (W8159, W11742);
not G9557 (W8160, I495);
not G9558 (W8161, W8162);
not G9559 (W8162, W11743);
not G9560 (W8163, I496);
not G9561 (W8164, W8165);
not G9562 (W8165, W11744);
not G9563 (W8166, I497);
not G9564 (W8167, W8169);
not G9565 (W8168, W11745);
not G9566 (W8169, W11746);
not G9567 (W8170, I498);
not G9568 (W8171, W8172);
not G9569 (W8172, W11747);
not G9570 (W8173, I499);
not G9571 (W8174, W8175);
not G9572 (W8175, W11748);
and G9573 (W8176, W11749, W11750);
and G9574 (W8177, I500, W11751);
and G9575 (W8178, W11752, W11753);
and G9576 (W8179, I501, W11754);
and G9577 (W8180, I502, W11755);
and G9578 (W8181, W11756, W11757);
and G9579 (W8182, I503, W11758);
and G9580 (W8183, W11759, W11760);
and G9581 (W8184, W11756, I500, W11761);
not G9582 (W8185, I504);
not G9583 (W8186, W8188);
not G9584 (W8187, W8242);
not G9585 (W8188, W11762);
not G9586 (W8189, I505);
not G9587 (W8190, W8192);
not G9588 (W8191, W8242);
not G9589 (W8192, W11763);
not G9590 (W8193, I506);
not G9591 (W8194, W8196);
not G9592 (W8195, W8242);
not G9593 (W8196, W11764);
not G9594 (W8197, I507);
not G9595 (W8198, W8200);
not G9596 (W8199, W8242);
not G9597 (W8200, W11765);
nand G9598 (W8201, W11766, W11767);
not G9599 (W8202, W8204);
not G9600 (W8203, I508);
not G9601 (W8204, W11768);
nand G9602 (W8205, W11769, W11770, W11771);
not G9603 (W8206, W8208);
not G9604 (W8207, I509);
not G9605 (W8208, W11772);
nand G9606 (W8209, W11773, W11774);
not G9607 (W8210, W8212);
not G9608 (W8211, I510);
not G9609 (W8212, W11775);
nand G9610 (W8213, W11776, W11777);
not G9611 (W8214, W8216);
not G9612 (W8215, I511);
not G9613 (W8216, W11778);
not G9614 (W8217, W8219);
not G9615 (W8218, I512);
not G9616 (W8219, W11779);
not G9617 (W8220, W8222);
not G9618 (W8221, I513);
not G9619 (W8222, W11780);
not G9620 (W8223, W8225);
not G9621 (W8224, I514);
not G9622 (W8225, W11781);
not G9623 (W8226, W8228);
not G9624 (W8227, I515);
not G9625 (W8228, W11782);
not G9626 (W8229, W8231);
not G9627 (W8230, I516);
not G9628 (W8231, W11783);
not G9629 (W8232, W8234);
not G9630 (W8233, I517);
not G9631 (W8234, W11784);
not G9632 (W8235, W8237);
not G9633 (W8236, I518);
not G9634 (W8237, W11785);
not G9635 (W8238, W8240);
not G9636 (W8239, I519);
not G9637 (W8240, W11786);
nand G9638 (W8241, W11787, W11788, W11789);
not G9639 (W8242, W11790);
not G9640 (W8243, W11791);
not G9641 (W8244, W11792);
nand G9642 (W8245, W11793, W11794);
not G9643 (W8246, W8248);
not G9644 (W8247, I520);
not G9645 (W8248, W11795);
nand G9646 (W8249, W11796, W11797, W11798);
not G9647 (W8250, W8252);
not G9648 (W8251, I521);
not G9649 (W8252, W11799);
nand G9650 (W8253, W11800, W11801);
not G9651 (W8254, W8256);
not G9652 (W8255, I522);
not G9653 (W8256, W11802);
nand G9654 (W8257, W11803, W11804);
not G9655 (W8258, W8260);
not G9656 (W8259, I523);
not G9657 (W8260, W11805);
not G9658 (W8261, W8263);
not G9659 (W8262, I524);
not G9660 (W8263, W11806);
not G9661 (W8264, W8266);
not G9662 (W8265, I525);
not G9663 (W8266, W11807);
not G9664 (W8267, W8269);
not G9665 (W8268, I526);
not G9666 (W8269, W11808);
not G9667 (W8270, W8272);
not G9668 (W8271, I527);
not G9669 (W8272, W11809);
not G9670 (W8273, W8275);
not G9671 (W8274, I528);
not G9672 (W8275, W11810);
not G9673 (W8276, W8278);
not G9674 (W8277, I529);
not G9675 (W8278, W11811);
not G9676 (W8279, W8281);
not G9677 (W8280, I530);
not G9678 (W8281, W11812);
not G9679 (W8282, W8284);
not G9680 (W8283, I531);
not G9681 (W8284, W11813);
nand G9682 (W8285, W11814, W11815, W11816);
not G9683 (W8286, W11817);
not G9684 (W8287, W11818);
nand G9685 (W8288, W11819, W11820);
not G9686 (W8289, W8291);
not G9687 (W8290, I532);
not G9688 (W8291, W11821);
nand G9689 (W8292, W11822, W11823, W11824);
not G9690 (W8293, W8295);
not G9691 (W8294, I533);
not G9692 (W8295, W11825);
nand G9693 (W8296, W11826, W11827);
not G9694 (W8297, W8299);
not G9695 (W8298, I534);
not G9696 (W8299, W11828);
nand G9697 (W8300, W11829, W11830);
not G9698 (W8301, W8303);
not G9699 (W8302, I535);
not G9700 (W8303, W11831);
not G9701 (W8304, W8306);
not G9702 (W8305, I536);
not G9703 (W8306, W11832);
not G9704 (W8307, W8309);
not G9705 (W8308, I537);
not G9706 (W8309, W11833);
not G9707 (W8310, W8312);
not G9708 (W8311, I538);
not G9709 (W8312, W11834);
not G9710 (W8313, W8315);
not G9711 (W8314, I539);
not G9712 (W8315, W11835);
not G9713 (W8316, W8318);
not G9714 (W8317, I540);
not G9715 (W8318, W11836);
not G9716 (W8319, W8321);
not G9717 (W8320, I541);
not G9718 (W8321, W11837);
not G9719 (W8322, W8324);
not G9720 (W8323, I542);
not G9721 (W8324, W11838);
not G9722 (W8325, W8327);
not G9723 (W8326, I543);
not G9724 (W8327, W11839);
nand G9725 (W8328, W11840, W11841, W11842);
not G9726 (W8329, W11843);
not G9727 (W8330, W11844);
nand G9728 (W8331, W11845, W11846);
not G9729 (W8332, W8334);
not G9730 (W8333, I544);
not G9731 (W8334, W11847);
nand G9732 (W8335, W11848, W11849, W11850);
not G9733 (W8336, W8338);
not G9734 (W8337, I545);
not G9735 (W8338, W11851);
nand G9736 (W8339, W11852, W11853);
not G9737 (W8340, W8342);
not G9738 (W8341, I546);
not G9739 (W8342, W11854);
nand G9740 (W8343, W11855, W11856);
not G9741 (W8344, W8346);
not G9742 (W8345, I547);
not G9743 (W8346, W11857);
not G9744 (W8347, W8349);
not G9745 (W8348, I548);
not G9746 (W8349, W11858);
not G9747 (W8350, W8352);
not G9748 (W8351, I549);
not G9749 (W8352, W11859);
not G9750 (W8353, W8355);
not G9751 (W8354, I550);
not G9752 (W8355, W11860);
not G9753 (W8356, W8358);
not G9754 (W8357, I551);
not G9755 (W8358, W11861);
not G9756 (W8359, W8361);
not G9757 (W8360, I552);
not G9758 (W8361, W11862);
not G9759 (W8362, W8364);
not G9760 (W8363, I553);
not G9761 (W8364, W11863);
not G9762 (W8365, W8367);
not G9763 (W8366, I554);
not G9764 (W8367, W11864);
not G9765 (W8368, W8370);
not G9766 (W8369, I555);
not G9767 (W8370, W11865);
nand G9768 (W8371, W11866, W11867, W11868);
not G9769 (W8372, W11869);
not G9770 (W8373, W11870);
and G9771 (W8374, I556, W11871);
and G9772 (W8375, W11872, W11873);
nor G9773 (W8376, W5847, W11874);
not G9774 (W8377, W8379);
nor G9775 (W8378, W11875, W11876);
not G9776 (W8379, W11877);
nor G9777 (W8380, W11878, W11879);
not G9778 (W8381, W8382);
not G9779 (W8382, W11880);
and G9780 (W8383, I557, W11881);
and G9781 (W8384, W11882, W11883);
and G9782 (W8385, W11884, W11885);
and G9783 (W8386, I558, W11886);
and G9784 (W8387, I559, W11887);
and G9785 (W8388, W11888, W11889);
and G9786 (W8389, W11890, W11891);
and G9787 (W8390, I560, W11892);
not G9788 (W8391, W11893);
not G9789 (W8392, W11894);
and G9790 (W8393, W11895, W11896);
and G9791 (W8394, W11897, W11898);
and G9792 (W8395, W11899, W11900);
and G9793 (W8396, W11901, W11902);
and G9794 (W8397, W11903, W11904);
and G9795 (W8398, W11905, W11906);
and G9796 (W8399, W11907, W11908);
and G9797 (W8400, W11909, W11910);
and G9798 (W8401, W11911, W11912);
and G9799 (W8402, W11913, W11914);
and G9800 (W8403, W11915, W11916);
and G9801 (W8404, W11917, W11918);
and G9802 (W8405, W11867, W11919);
and G9803 (W8406, W11920, W11921);
and G9804 (W8407, W11922, W11923);
and G9805 (W8408, W11924, W11925);
and G9806 (W8409, W11926, W11927);
and G9807 (W8410, W11928, W11929);
and G9808 (W8411, W11930, W11931);
not G9809 (W8412, W11932);
not G9810 (W8413, W8415);
not G9811 (W8414, I561);
not G9812 (W8415, W11933);
not G9813 (W8416, W8418);
not G9814 (W8417, I562);
not G9815 (W8418, W11934);
not G9816 (W8419, W8421);
not G9817 (W8420, I563);
not G9818 (W8421, W11935);
not G9819 (W8422, W11936);
not G9820 (W8423, W8425);
not G9821 (W8424, I564);
not G9822 (W8425, W11937);
not G9823 (W8426, W8428);
not G9824 (W8427, I565);
not G9825 (W8428, W11938);
not G9826 (W8429, W8431);
not G9827 (W8430, I566);
not G9828 (W8431, W11939);
not G9829 (W8432, W11940);
not G9830 (W8433, W8435);
not G9831 (W8434, I567);
not G9832 (W8435, W11941);
not G9833 (W8436, W8438);
not G9834 (W8437, I568);
not G9835 (W8438, W11942);
not G9836 (W8439, W8441);
not G9837 (W8440, I569);
not G9838 (W8441, W11943);
not G9839 (W8442, W11944);
not G9840 (W8443, W8445);
not G9841 (W8444, I570);
not G9842 (W8445, W11945);
not G9843 (W8446, W8448);
not G9844 (W8447, I571);
not G9845 (W8448, W11946);
not G9846 (W8449, W8451);
not G9847 (W8450, I572);
not G9848 (W8451, W11947);
not G9849 (W8452, W8454);
not G9850 (W8453, I573);
not G9851 (W8454, W11948);
not G9852 (W8455, W8457);
not G9853 (W8456, I574);
not G9854 (W8457, W11949);
not G9855 (W8458, W8460);
not G9856 (W8459, I575);
not G9857 (W8460, W11950);
not G9858 (W8461, W8463);
not G9859 (W8462, I576);
not G9860 (W8463, W11951);
not G9861 (W8464, W8466);
not G9862 (W8465, I577);
not G9863 (W8466, W11952);
not G9864 (W8467, W8469);
not G9865 (W8468, I578);
not G9866 (W8469, W11953);
not G9867 (W8470, W8472);
not G9868 (W8471, I579);
not G9869 (W8472, W11954);
not G9870 (W8473, W8475);
not G9871 (W8474, I580);
not G9872 (W8475, W11955);
not G9873 (W8476, W8478);
not G9874 (W8477, I581);
not G9875 (W8478, W11956);
not G9876 (W8479, W8481);
not G9877 (W8480, I582);
not G9878 (W8481, W11957);
not G9879 (W8482, W8484);
not G9880 (W8483, I583);
not G9881 (W8484, W11958);
not G9882 (W8485, W8487);
not G9883 (W8486, I584);
not G9884 (W8487, W11959);
not G9885 (W8488, W8490);
not G9886 (W8489, I585);
not G9887 (W8490, W11960);
not G9888 (W8491, W8493);
not G9889 (W8492, I586);
not G9890 (W8493, W11961);
not G9891 (W8494, W8496);
not G9892 (W8495, I587);
not G9893 (W8496, W11962);
not G9894 (W8497, W8499);
not G9895 (W8498, I588);
not G9896 (W8499, W11963);
not G9897 (W8500, W8502);
not G9898 (W8501, I589);
not G9899 (W8502, W11964);
not G9900 (W8503, W8505);
not G9901 (W8504, I590);
not G9902 (W8505, W11965);
not G9903 (W8506, W8508);
not G9904 (W8507, I591);
not G9905 (W8508, W11966);
not G9906 (W8509, W8511);
not G9907 (W8510, I592);
not G9908 (W8511, W11967);
not G9909 (W8512, W8514);
not G9910 (W8513, I593);
not G9911 (W8514, W11968);
not G9912 (W8515, W8517);
not G9913 (W8516, I594);
not G9914 (W8517, W11969);
not G9915 (W8518, W8520);
not G9916 (W8519, I595);
not G9917 (W8520, W11970);
not G9918 (W8521, W8523);
not G9919 (W8522, I596);
not G9920 (W8523, W11971);
not G9921 (W8524, W8526);
not G9922 (W8525, I597);
not G9923 (W8526, W11972);
not G9924 (W8527, W8529);
not G9925 (W8528, I598);
not G9926 (W8529, W11973);
not G9927 (W8530, W8532);
not G9928 (W8531, I599);
not G9929 (W8532, W11974);
not G9930 (W8533, W8535);
not G9931 (W8534, I600);
not G9932 (W8535, W11975);
not G9933 (W8536, W8538);
not G9934 (W8537, I601);
not G9935 (W8538, W11976);
not G9936 (W8539, W8541);
not G9937 (W8540, I602);
not G9938 (W8541, W11977);
and G9939 (W8542, I260, W11978);
and G9940 (W8543, W11979, W11980);
not G9941 (W8544, W11981);
and G9942 (W8545, W11982, W11983);
and G9943 (W8546, I261, W11984);
and G9944 (W8547, I262, W11985);
and G9945 (W8548, W11986, W11987);
and G9946 (W8549, W11988, W11989);
and G9947 (W8550, I263, W11990);
and G9948 (W8551, I264, W11991);
and G9949 (W8552, W11992, W11993);
and G9950 (W8553, W11994, W11995);
and G9951 (W8554, I265, W11996);
and G9952 (W8555, I266, W11997);
and G9953 (W8556, W11998, W11999);
and G9954 (W8557, W12000, W12001);
and G9955 (W8558, I267, W12002);
and G9956 (W8559, I268, W12003);
and G9957 (W8560, W12004, W12005);
and G9958 (W8561, W12006, W12007);
and G9959 (W8562, I269, W12008);
not G9960 (W8563, I603);
not G9961 (W8564, W8566);
not G9962 (W8565, I604);
not G9963 (W8566, W12009);
nor G9964 (W8567, W12010, W12011);
not G9965 (W8568, W8570);
not G9966 (W8569, I605);
not G9967 (W8570, W12012);
nor G9968 (W8571, W12013, W12014);
not G9969 (W8572, W8574);
not G9970 (W8573, I606);
not G9971 (W8574, W12015);
nor G9972 (W8575, W12016, W12017);
not G9973 (W8576, W8578);
not G9974 (W8577, I607);
not G9975 (W8578, W12018);
nor G9976 (W8579, W12019, W12020);
not G9977 (W8580, W8582);
not G9978 (W8581, I608);
not G9979 (W8582, W12021);
nor G9980 (W8583, W12022, W12023);
not G9981 (W8584, W8586);
not G9982 (W8585, I609);
not G9983 (W8586, W12024);
not G9984 (W8587, I610);
not G9985 (W8588, W8590);
not G9986 (W8589, W12025);
not G9987 (W8590, W12026);
not G9988 (W8591, I611);
not G9989 (W8592, W8593);
not G9990 (W8593, W12027);
not G9991 (W8594, I612);
not G9992 (W8595, W8596);
not G9993 (W8596, W12028);
and G9994 (W8597, W8696, W8369);
and G9995 (W8598, W8697, W8366);
and G9996 (W8599, W8698, W8345);
and G9997 (W8600, W8696, W8363);
and G9998 (W8601, W8697, W8360);
and G9999 (W8602, W8698, W8341);
and G10000 (W8603, W8696, W8357);
and G10001 (W8604, W8697, W8354);
and G10002 (W8605, W8698, W8337);
and G10003 (W8606, W8696, W8351);
and G10004 (W8607, W8697, W8348);
and G10005 (W8608, W8698, W8333);
not G10006 (W8609, I613);
not G10007 (W8610, W8612);
not G10008 (W8611, W12029);
not G10009 (W8612, W12030);
not G10010 (W8613, I614);
not G10011 (W8614, W8615);
not G10012 (W8615, W12031);
not G10013 (W8616, I615);
not G10014 (W8617, W8618);
not G10015 (W8618, W12032);
not G10016 (W8619, I616);
not G10017 (W8620, W8622);
not G10018 (W8621, W12033);
not G10019 (W8622, W12034);
not G10020 (W8623, I617);
not G10021 (W8624, W8625);
not G10022 (W8625, W12035);
not G10023 (W8626, I618);
not G10024 (W8627, W8628);
not G10025 (W8628, W12036);
nor G10026 (W8629, W12037, W12038);
not G10027 (W8630, W8632);
not G10028 (W8631, I619);
not G10029 (W8632, W12039);
not G10030 (W8633, I620);
not G10031 (W8634, W8636);
not G10032 (W8635, W12040);
not G10033 (W8636, W12041);
not G10034 (W8637, I621);
not G10035 (W8638, W8639);
not G10036 (W8639, W12042);
not G10037 (W8640, I622);
not G10038 (W8641, W8642);
not G10039 (W8642, W12043);
not G10040 (W8643, I270);
not G10041 (W8644, W8646);
not G10042 (W8645, W12044);
not G10043 (W8646, W12045);
not G10044 (W8647, I271);
not G10045 (W8648, W8649);
not G10046 (W8649, W12046);
not G10047 (W8650, I272);
not G10048 (W8651, W8652);
not G10049 (W8652, W12047);
nor G10050 (W8653, W12048, W12049, W12050);
not G10051 (W8654, I623);
not G10052 (W8655, W8657);
not G10053 (W8656, W12051);
not G10054 (W8657, W12052);
not G10055 (W8658, I624);
not G10056 (W8659, W8660);
not G10057 (W8660, W12053);
not G10058 (W8661, I625);
not G10059 (W8662, W8663);
not G10060 (W8663, W12054);
nor G10061 (W8664, W12055, W12056, W12057);
not G10062 (W8665, I626);
not G10063 (W8666, W8668);
not G10064 (W8667, W12058);
not G10065 (W8668, W12059);
not G10066 (W8669, I627);
not G10067 (W8670, W8671);
not G10068 (W8671, W12060);
not G10069 (W8672, I628);
not G10070 (W8673, W8674);
not G10071 (W8674, W12061);
not G10072 (W8675, I273);
not G10073 (W8676, W8678);
not G10074 (W8677, W12062);
not G10075 (W8678, W12063);
not G10076 (W8679, I274);
not G10077 (W8680, W8681);
not G10078 (W8681, W12064);
not G10079 (W8682, I275);
not G10080 (W8683, W8684);
not G10081 (W8684, W12065);
nor G10082 (W8685, W12066, W12067, W12068);
not G10083 (W8686, I629);
not G10084 (W8687, W8689);
not G10085 (W8688, W12069);
not G10086 (W8689, W12070);
not G10087 (W8690, I630);
not G10088 (W8691, W8692);
not G10089 (W8692, W12071);
not G10090 (W8693, I631);
not G10091 (W8694, W8695);
not G10092 (W8695, W12072);
not G10093 (W8696, W12073);
not G10094 (W8697, W12074);
not G10095 (W8698, W12075);
not G10096 (W8699, I604);
not G10097 (W8700, W8702);
not G10098 (W8701, I632);
not G10099 (W8702, W12076);
not G10100 (W8703, W8704);
not G10101 (W8704, W12077);
nor G10102 (W8705, W12078, W12079);
not G10103 (W8706, W8707);
not G10104 (W8707, W12080);
nor G10105 (W8708, W12081, W12082);
not G10106 (W8709, W8711);
not G10107 (W8710, I633);
not G10108 (W8711, W12083);
nor G10109 (W8712, W12084, W12085);
not G10110 (W8713, W8715);
not G10111 (W8714, I634);
not G10112 (W8715, W12086);
nor G10113 (W8716, W12087, W12088);
not G10114 (W8717, W8719);
not G10115 (W8718, I635);
not G10116 (W8719, W12089);
nor G10117 (W8720, W12090, W12091);
not G10118 (W8721, W8723);
not G10119 (W8722, I636);
not G10120 (W8723, W12092);
nor G10121 (W8724, W12093, W12094);
not G10122 (W8725, W8727);
not G10123 (W8726, I637);
not G10124 (W8727, W12095);
nor G10125 (W8728, W12096, W12097);
not G10126 (W8729, I638);
not G10127 (W8730, I639);
not G10128 (W8731, I640);
not G10129 (W8732, I641);
not G10130 (W8733, I642);
not G10131 (W8734, I643);
not G10132 (W8735, I644);
not G10133 (W8736, I645);
not G10134 (W8737, I646);
and G10135 (W8738, W12098, W12099);
not G10136 (W8739, W8741);
not G10137 (W8740, I647);
not G10138 (W8741, W12100);
not G10139 (W8742, W8744);
not G10140 (W8743, I648);
not G10141 (W8744, W12101);
not G10142 (W8745, W8747);
not G10143 (W8746, I649);
not G10144 (W8747, W12102);
not G10145 (W8748, I650);
not G10146 (W8749, W8751);
not G10147 (W8750, W12103);
not G10148 (W8751, W12104);
not G10149 (W8752, I651);
not G10150 (W8753, W8754);
not G10151 (W8754, W12105);
not G10152 (W8755, I652);
not G10153 (W8756, W8757);
not G10154 (W8757, W12106);
not G10155 (W8758, I653);
not G10156 (W8759, W8761);
not G10157 (W8760, W12107);
not G10158 (W8761, W12108);
not G10159 (W8762, I654);
not G10160 (W8763, W8764);
not G10161 (W8764, W12109);
not G10162 (W8765, I655);
not G10163 (W8766, W8767);
not G10164 (W8767, W12110);
not G10165 (W8768, I656);
not G10166 (W8769, W8771);
not G10167 (W8770, W12111);
not G10168 (W8771, W12112);
not G10169 (W8772, I657);
not G10170 (W8773, W8774);
not G10171 (W8774, W12113);
not G10172 (W8775, I658);
not G10173 (W8776, W8777);
not G10174 (W8777, W12114);
not G10175 (W8778, I659);
not G10176 (W8779, W8781);
not G10177 (W8780, W12115);
not G10178 (W8781, W12116);
not G10179 (W8782, I660);
not G10180 (W8783, W8784);
not G10181 (W8784, W12117);
not G10182 (W8785, I661);
not G10183 (W8786, W8787);
not G10184 (W8787, W12118);
not G10185 (W8788, I662);
not G10186 (W8789, W8791);
not G10187 (W8790, W12119);
not G10188 (W8791, W12120);
not G10189 (W8792, I663);
not G10190 (W8793, W8794);
not G10191 (W8794, W12121);
not G10192 (W8795, I664);
not G10193 (W8796, W8797);
not G10194 (W8797, W12122);
not G10195 (W8798, I665);
not G10196 (W8799, W8801);
not G10197 (W8800, W12123);
not G10198 (W8801, W12124);
not G10199 (W8802, I666);
not G10200 (W8803, W8804);
not G10201 (W8804, W12125);
not G10202 (W8805, I667);
not G10203 (W8806, W8807);
not G10204 (W8807, W12126);
not G10205 (W8808, I668);
not G10206 (W8809, W8811);
not G10207 (W8810, W12127);
not G10208 (W8811, W12128);
not G10209 (W8812, I669);
not G10210 (W8813, W8814);
not G10211 (W8814, W12129);
not G10212 (W8815, I670);
not G10213 (W8816, W8817);
not G10214 (W8817, W12130);
not G10215 (W8818, I671);
not G10216 (W8819, W8821);
not G10217 (W8820, W12131);
not G10218 (W8821, W12132);
not G10219 (W8822, I672);
not G10220 (W8823, W8824);
not G10221 (W8824, W12133);
not G10222 (W8825, I673);
not G10223 (W8826, W8827);
not G10224 (W8827, W12134);
not G10225 (W8828, I674);
not G10226 (W8829, W8831);
not G10227 (W8830, W12135);
not G10228 (W8831, W12136);
not G10229 (W8832, I675);
not G10230 (W8833, W8834);
not G10231 (W8834, W12137);
not G10232 (W8835, I676);
not G10233 (W8836, W8837);
not G10234 (W8837, W12138);
not G10235 (W8838, I677);
not G10236 (W8839, W8841);
not G10237 (W8840, W12139);
not G10238 (W8841, W12140);
not G10239 (W8842, I678);
not G10240 (W8843, W8844);
not G10241 (W8844, W12141);
not G10242 (W8845, I679);
not G10243 (W8846, W8847);
not G10244 (W8847, W12142);
not G10245 (W8848, I680);
not G10246 (W8849, W8851);
not G10247 (W8850, W12143);
not G10248 (W8851, W12144);
not G10249 (W8852, I681);
not G10250 (W8853, W8854);
not G10251 (W8854, W12145);
not G10252 (W8855, I682);
not G10253 (W8856, W8857);
not G10254 (W8857, W12146);
not G10255 (W8858, I683);
not G10256 (W8859, W8861);
not G10257 (W8860, W12147);
not G10258 (W8861, W12148);
not G10259 (W8862, I684);
not G10260 (W8863, W8864);
not G10261 (W8864, W12149);
not G10262 (W8865, I685);
not G10263 (W8866, W8867);
not G10264 (W8867, W12150);
not G10265 (W8868, I686);
not G10266 (W8869, W8871);
not G10267 (W8870, W12151);
not G10268 (W8871, W12152);
not G10269 (W8872, I687);
not G10270 (W8873, W8874);
not G10271 (W8874, W12153);
not G10272 (W8875, I688);
not G10273 (W8876, W8877);
not G10274 (W8877, W12154);
nor G10275 (W8878, W12155, W12156);
not G10276 (W8879, W8881);
not G10277 (W8880, I689);
not G10278 (W8881, W12157);
not G10279 (W8882, W8884);
not G10280 (W8883, I690);
not G10281 (W8884, W12158);
not G10282 (W8885, W8887);
not G10283 (W8886, I691);
not G10284 (W8887, W12159);
not G10285 (W8888, W12160);
nor G10286 (W8889, W12161, W12162);
nand G10287 (W8890, W12163, W12164);
not G10288 (W8891, W8893);
not G10289 (W8892, I293);
not G10290 (W8893, W12165);
nand G10291 (W8894, W12166, W12167, W12168);
not G10292 (W8895, W8897);
not G10293 (W8896, I290);
not G10294 (W8897, W12169);
nand G10295 (W8898, W12170, W12171);
not G10296 (W8899, W8901);
not G10297 (W8900, I287);
not G10298 (W8901, W12172);
nand G10299 (W8902, W12173, W12174);
not G10300 (W8903, W8905);
not G10301 (W8904, I284);
not G10302 (W8905, W12175);
not G10303 (W8906, W8908);
not G10304 (W8907, I294);
not G10305 (W8908, W12176);
not G10306 (W8909, W8911);
not G10307 (W8910, I295);
not G10308 (W8911, W12177);
not G10309 (W8912, W8914);
not G10310 (W8913, I291);
not G10311 (W8914, W12178);
not G10312 (W8915, W8917);
not G10313 (W8916, I292);
not G10314 (W8917, W12179);
not G10315 (W8918, W8920);
not G10316 (W8919, I288);
not G10317 (W8920, W12180);
not G10318 (W8921, W8923);
not G10319 (W8922, I289);
not G10320 (W8923, W12181);
not G10321 (W8924, W8926);
not G10322 (W8925, I285);
not G10323 (W8926, W12182);
not G10324 (W8927, W8929);
not G10325 (W8928, I286);
not G10326 (W8929, W12183);
not G10327 (W8930, I692);
not G10328 (W8931, W8933);
not G10329 (W8932, W12184);
not G10330 (W8933, W12185);
not G10331 (W8934, I693);
not G10332 (W8935, W8936);
not G10333 (W8936, W12186);
not G10334 (W8937, I694);
not G10335 (W8938, W8939);
not G10336 (W8939, W12187);
nor G10337 (W8940, W12188, W12189, W12190);
not G10338 (W8941, W8943);
not G10339 (W8942, I695);
not G10340 (W8943, W12191);
not G10341 (W8944, W8946);
not G10342 (W8945, I696);
not G10343 (W8946, W12192);
not G10344 (W8947, W8949);
not G10345 (W8948, I697);
not G10346 (W8949, W12193);
not G10347 (W8950, I698);
not G10348 (W8951, W8953);
not G10349 (W8952, W12194);
not G10350 (W8953, W12195);
not G10351 (W8954, I699);
not G10352 (W8955, W8956);
not G10353 (W8956, W12196);
not G10354 (W8957, I700);
not G10355 (W8958, W8959);
not G10356 (W8959, W12197);
not G10357 (W8960, I701);
not G10358 (W8961, W8963);
not G10359 (W8962, W12198);
not G10360 (W8963, W12199);
not G10361 (W8964, I702);
not G10362 (W8965, W8966);
not G10363 (W8966, W12200);
not G10364 (W8967, I703);
not G10365 (W8968, W8969);
not G10366 (W8969, W12201);
not G10367 (W8970, I704);
not G10368 (W8971, W8973);
not G10369 (W8972, W12202);
not G10370 (W8973, W12203);
not G10371 (W8974, I705);
not G10372 (W8975, W8976);
not G10373 (W8976, W12204);
not G10374 (W8977, I706);
not G10375 (W8978, W8979);
not G10376 (W8979, W12205);
not G10377 (W8980, W12206);
not G10378 (W8981, W8983);
not G10379 (W8982, I707);
not G10380 (W8983, W12207);
not G10381 (W8984, W8986);
not G10382 (W8985, I708);
not G10383 (W8986, W12208);
not G10384 (W8987, W8989);
not G10385 (W8988, I709);
not G10386 (W8989, W12209);
and G10387 (W8990, W12210, I701);
and G10388 (W8991, W12211, I702);
and G10389 (W8992, W12212, I703);
and G10390 (W8993, W12210, W8928);
and G10391 (W8994, W12211, W8925);
and G10392 (W8995, W12212, W8904);
and G10393 (W8996, W12210, W8922);
and G10394 (W8997, W12211, W8919);
and G10395 (W8998, W12212, W8900);
and G10396 (W8999, W12210, W8916);
and G10397 (W9000, W12211, W8913);
and G10398 (W9001, W12212, W8896);
and G10399 (W9002, W12210, W8910);
and G10400 (W9003, W12211, W8907);
and G10401 (W9004, W12212, W8892);
not G10402 (W9005, W12213);
not G10403 (W9006, W9008);
not G10404 (W9007, I710);
not G10405 (W9008, W12214);
not G10406 (W9009, W12215);
not G10407 (W9010, W9012);
not G10408 (W9011, I711);
not G10409 (W9012, W12216);
not G10410 (W9013, W12217);
not G10411 (W9014, W9016);
not G10412 (W9015, I712);
not G10413 (W9016, W12218);
not G10414 (W9017, W12219);
not G10415 (W9018, W9020);
not G10416 (W9019, I713);
not G10417 (W9020, W12220);
not G10418 (W9021, W12221);
not G10419 (W9022, W9024);
not G10420 (W9023, I714);
not G10421 (W9024, W12222);
not G10422 (W9025, W12223);
not G10423 (W9026, W9028);
not G10424 (W9027, I715);
not G10425 (W9028, W12224);
not G10426 (W9029, W12225);
not G10427 (W9030, W9032);
not G10428 (W9031, I716);
not G10429 (W9032, W12226);
not G10430 (W9033, W12227);
not G10431 (W9034, W9036);
not G10432 (W9035, I717);
not G10433 (W9036, W12228);
not G10434 (W9037, W12229);
not G10435 (W9038, W9040);
not G10436 (W9039, I718);
not G10437 (W9040, W12230);
not G10438 (W9041, W12231);
not G10439 (W9042, W9044);
not G10440 (W9043, I719);
not G10441 (W9044, W12232);
not G10442 (W9045, W9047);
not G10443 (W9046, I720);
not G10444 (W9047, W12233);
not G10445 (W9048, W9050);
not G10446 (W9049, I721);
not G10447 (W9050, W12234);
not G10448 (W9051, W9053);
not G10449 (W9052, I722);
not G10450 (W9053, W12235);
not G10451 (W9054, W9056);
not G10452 (W9055, I723);
not G10453 (W9056, W12236);
not G10454 (W9057, W9059);
not G10455 (W9058, I724);
not G10456 (W9059, W12237);
not G10457 (W9060, W9062);
not G10458 (W9061, I725);
not G10459 (W9062, W12238);
not G10460 (W9063, W9065);
not G10461 (W9064, I726);
not G10462 (W9065, W12239);
not G10463 (W9066, W9068);
not G10464 (W9067, I727);
not G10465 (W9068, W12240);
not G10466 (W9069, W9071);
not G10467 (W9070, I728);
not G10468 (W9071, W12241);
not G10469 (W9072, W9074);
not G10470 (W9073, I729);
not G10471 (W9074, W12242);
not G10472 (W9075, W9077);
not G10473 (W9076, I730);
not G10474 (W9077, W12243);
not G10475 (W9078, W9080);
not G10476 (W9079, I731);
not G10477 (W9080, W12244);
not G10478 (W9081, W9083);
not G10479 (W9082, I732);
not G10480 (W9083, W12245);
not G10481 (W9084, W9086);
not G10482 (W9085, I733);
not G10483 (W9086, W12246);
not G10484 (W9087, W9089);
not G10485 (W9088, I734);
not G10486 (W9089, W12247);
not G10487 (W9090, W9092);
not G10488 (W9091, I735);
not G10489 (W9092, W12248);
not G10490 (W9093, W9095);
not G10491 (W9094, I736);
not G10492 (W9095, W12249);
not G10493 (W9096, W9098);
not G10494 (W9097, I737);
not G10495 (W9098, W12250);
not G10496 (W9099, W9101);
not G10497 (W9100, I738);
not G10498 (W9101, W12251);
not G10499 (W9102, W9104);
not G10500 (W9103, I739);
not G10501 (W9104, W12252);
and G10502 (W9105, I740, W12253);
and G10503 (W9106, W12254, W12255);
not G10504 (W9107, W12256);
not G10505 (W9108, W12257);
not G10506 (W9109, W12258);
and G10507 (W9110, W12259, W12260);
and G10508 (W9111, I741, W12261);
and G10509 (W9112, I742, W12262);
and G10510 (W9113, W12263, W12264);
and G10511 (W9114, W12265, W12266);
and G10512 (W9115, I743, W12267);
and G10513 (W9116, I744, W12268);
and G10514 (W9117, W12269, W12270);
and G10515 (W9118, W12271, W12272);
and G10516 (W9119, I745, W12273);
and G10517 (W9120, I746, W12274);
and G10518 (W9121, W12275, W12276);
and G10519 (W9122, W12277, W12278);
and G10520 (W9123, I747, W12279);
and G10521 (W9124, I748, W12280);
and G10522 (W9125, W12281, W12282);
and G10523 (W9126, W12283, W12284);
and G10524 (W9127, I749, W12285);
and G10525 (W9128, W12286, W12287);
not G10526 (W9129, W9131);
not G10527 (W9130, I750);
not G10528 (W9131, W12288);
not G10529 (W9132, W9134);
not G10530 (W9133, I751);
not G10531 (W9134, W12289);
not G10532 (W9135, W9137);
not G10533 (W9136, I752);
not G10534 (W9137, W12290);
not G10535 (W9138, W9140);
not G10536 (W9139, I753);
not G10537 (W9140, W12291);
not G10538 (W9141, W9143);
not G10539 (W9142, I754);
not G10540 (W9143, W12292);
not G10541 (W9144, W9146);
not G10542 (W9145, I755);
not G10543 (W9146, W12293);
not G10544 (W9147, W9149);
not G10545 (W9148, I756);
not G10546 (W9149, W12294);
not G10547 (W9150, W9152);
not G10548 (W9151, I757);
not G10549 (W9152, W12295);
not G10550 (W9153, W9155);
not G10551 (W9154, I758);
not G10552 (W9155, W12296);
nand G10553 (W9156, W9013, W9025, W12297);
not G10554 (W9157, W9159);
not G10555 (W9158, I759);
not G10556 (W9159, W12298);
not G10557 (W9160, W9162);
not G10558 (W9161, I760);
not G10559 (W9162, W12299);
not G10560 (W9163, W9165);
not G10561 (W9164, I761);
not G10562 (W9165, W12300);
and G10563 (W9166, W12301, W12302);
and G10564 (W9167, W12303, W12304);
and G10565 (W9168, W12305, W12306);
and G10566 (W9169, W12307, W12308);
and G10567 (W9170, W12309, W12310);
and G10568 (W9171, W12311, W12312);
and G10569 (W9172, W12313, W12314);
and G10570 (W9173, W12315, W12316);
and G10571 (W9174, W12317, W12318);
and G10572 (W9175, W12319, W12320);
and G10573 (W9176, W12321, W12322);
and G10574 (W9177, W12323, W12324);
and G10575 (W9178, W11841, W12325);
and G10576 (W9179, W12326, W12327);
and G10577 (W9180, W12328, W12329);
and G10578 (W9181, W12330, W12331);
and G10579 (W9182, W12332, W12333);
and G10580 (W9183, W12334, W12335);
and G10581 (W9184, W12336, W12337);
not G10582 (W9185, W12338);
not G10583 (W9186, W9188);
not G10584 (W9187, I762);
not G10585 (W9188, W12339);
not G10586 (W9189, W9191);
not G10587 (W9190, I763);
not G10588 (W9191, W12340);
not G10589 (W9192, W9194);
not G10590 (W9193, I764);
not G10591 (W9194, W12341);
not G10592 (W9195, W12342);
not G10593 (W9196, W9198);
not G10594 (W9197, I765);
not G10595 (W9198, W12343);
not G10596 (W9199, W9201);
not G10597 (W9200, I766);
not G10598 (W9201, W12344);
not G10599 (W9202, W9204);
not G10600 (W9203, I767);
not G10601 (W9204, W12345);
not G10602 (W9205, W12346);
not G10603 (W9206, W9208);
not G10604 (W9207, I768);
not G10605 (W9208, W12347);
not G10606 (W9209, W9211);
not G10607 (W9210, I769);
not G10608 (W9211, W12348);
not G10609 (W9212, W9214);
not G10610 (W9213, I770);
not G10611 (W9214, W12349);
not G10612 (W9215, W12350);
not G10613 (W9216, W9218);
not G10614 (W9217, I771);
not G10615 (W9218, W12351);
not G10616 (W9219, W9221);
not G10617 (W9220, I772);
not G10618 (W9221, W12352);
not G10619 (W9222, W9224);
not G10620 (W9223, I773);
not G10621 (W9224, W12353);
not G10622 (W9225, W9227);
not G10623 (W9226, I774);
not G10624 (W9227, W12354);
not G10625 (W9228, W9230);
not G10626 (W9229, I775);
not G10627 (W9230, W12355);
not G10628 (W9231, W9233);
not G10629 (W9232, I776);
not G10630 (W9233, W12356);
not G10631 (W9234, W9236);
not G10632 (W9235, I777);
not G10633 (W9236, W12357);
not G10634 (W9237, W9239);
not G10635 (W9238, I778);
not G10636 (W9239, W12358);
not G10637 (W9240, W9242);
not G10638 (W9241, I779);
not G10639 (W9242, W12359);
not G10640 (W9243, W9245);
not G10641 (W9244, I780);
not G10642 (W9245, W12360);
not G10643 (W9246, W9248);
not G10644 (W9247, I781);
not G10645 (W9248, W12361);
not G10646 (W9249, W9251);
not G10647 (W9250, I782);
not G10648 (W9251, W12362);
not G10649 (W9252, W9254);
not G10650 (W9253, I783);
not G10651 (W9254, W12363);
not G10652 (W9255, W9257);
not G10653 (W9256, I784);
not G10654 (W9257, W12364);
not G10655 (W9258, W9260);
not G10656 (W9259, I785);
not G10657 (W9260, W12365);
not G10658 (W9261, W9263);
not G10659 (W9262, I786);
not G10660 (W9263, W12366);
not G10661 (W9264, W9266);
not G10662 (W9265, I787);
not G10663 (W9266, W12367);
not G10664 (W9267, W9269);
not G10665 (W9268, I788);
not G10666 (W9269, W12368);
not G10667 (W9270, W9272);
not G10668 (W9271, I789);
not G10669 (W9272, W12369);
not G10670 (W9273, W9275);
not G10671 (W9274, I790);
not G10672 (W9275, W12370);
not G10673 (W9276, W9278);
not G10674 (W9277, I791);
not G10675 (W9278, W12371);
not G10676 (W9279, W9281);
not G10677 (W9280, I792);
not G10678 (W9281, W12372);
not G10679 (W9282, W9284);
not G10680 (W9283, I793);
not G10681 (W9284, W12373);
not G10682 (W9285, W9287);
not G10683 (W9286, I794);
not G10684 (W9287, W12374);
not G10685 (W9288, W9290);
not G10686 (W9289, I795);
not G10687 (W9290, W12375);
not G10688 (W9291, W9293);
not G10689 (W9292, I796);
not G10690 (W9293, W12376);
not G10691 (W9294, W9296);
not G10692 (W9295, I797);
not G10693 (W9296, W12377);
not G10694 (W9297, W9299);
not G10695 (W9298, I798);
not G10696 (W9299, W12378);
not G10697 (W9300, W9302);
not G10698 (W9301, I799);
not G10699 (W9302, W12379);
not G10700 (W9303, W9305);
not G10701 (W9304, I800);
not G10702 (W9305, W12380);
not G10703 (W9306, W9308);
not G10704 (W9307, I801);
not G10705 (W9308, W12381);
not G10706 (W9309, W9311);
not G10707 (W9310, I802);
not G10708 (W9311, W12382);
not G10709 (W9312, W9314);
not G10710 (W9313, I803);
not G10711 (W9314, W12383);
and G10712 (W9315, I296, W12384);
and G10713 (W9316, W12385, W12386);
not G10714 (W9317, W12387);
and G10715 (W9318, W12388, W12389);
and G10716 (W9319, I297, W12390);
and G10717 (W9320, I298, W12391);
and G10718 (W9321, W12392, W12393);
and G10719 (W9322, W12394, W12395);
and G10720 (W9323, I299, W12396);
and G10721 (W9324, I300, W12397);
and G10722 (W9325, W12398, W12399);
and G10723 (W9326, W12400, W12401);
and G10724 (W9327, I301, W12402);
and G10725 (W9328, I302, W12403);
and G10726 (W9329, W12404, W12405);
and G10727 (W9330, W12406, W12407);
and G10728 (W9331, I303, W12408);
and G10729 (W9332, I304, W12409);
and G10730 (W9333, W12410, W12411);
and G10731 (W9334, W12412, W12413);
and G10732 (W9335, I305, W12414);
not G10733 (W9336, I804);
not G10734 (W9337, W9339);
not G10735 (W9338, I805);
not G10736 (W9339, W12415);
nor G10737 (W9340, W12416, W12417);
not G10738 (W9341, W9343);
not G10739 (W9342, I806);
not G10740 (W9343, W12418);
nor G10741 (W9344, W12419, W12420);
not G10742 (W9345, W9347);
not G10743 (W9346, I807);
not G10744 (W9347, W12421);
nor G10745 (W9348, W12422, W12423);
not G10746 (W9349, W9351);
not G10747 (W9350, I808);
not G10748 (W9351, W12424);
nor G10749 (W9352, W12425, W12426);
not G10750 (W9353, W9355);
not G10751 (W9354, I809);
not G10752 (W9355, W12427);
nor G10753 (W9356, W12428, W12429);
not G10754 (W9357, W9359);
not G10755 (W9358, I810);
not G10756 (W9359, W12430);
not G10757 (W9360, I811);
not G10758 (W9361, W9363);
not G10759 (W9362, W12431);
not G10760 (W9363, W12432);
not G10761 (W9364, I812);
not G10762 (W9365, W9366);
not G10763 (W9366, W12433);
not G10764 (W9367, I813);
not G10765 (W9368, W9369);
not G10766 (W9369, W12434);
and G10767 (W9370, W9469, W8326);
and G10768 (W9371, W9470, W8323);
and G10769 (W9372, W9471, W8302);
and G10770 (W9373, W9469, W8320);
and G10771 (W9374, W9470, W8317);
and G10772 (W9375, W9471, W8298);
and G10773 (W9376, W9469, W8314);
and G10774 (W9377, W9470, W8311);
and G10775 (W9378, W9471, W8294);
and G10776 (W9379, W9469, W8308);
and G10777 (W9380, W9470, W8305);
and G10778 (W9381, W9471, W8290);
not G10779 (W9382, I814);
not G10780 (W9383, W9385);
not G10781 (W9384, W12435);
not G10782 (W9385, W12436);
not G10783 (W9386, I815);
not G10784 (W9387, W9388);
not G10785 (W9388, W12437);
not G10786 (W9389, I816);
not G10787 (W9390, W9391);
not G10788 (W9391, W12438);
not G10789 (W9392, I817);
not G10790 (W9393, W9395);
not G10791 (W9394, W12439);
not G10792 (W9395, W12440);
not G10793 (W9396, I818);
not G10794 (W9397, W9398);
not G10795 (W9398, W12441);
not G10796 (W9399, I819);
not G10797 (W9400, W9401);
not G10798 (W9401, W12442);
nor G10799 (W9402, W12443, W12444);
not G10800 (W9403, W9405);
not G10801 (W9404, I820);
not G10802 (W9405, W12445);
not G10803 (W9406, I821);
not G10804 (W9407, W9409);
not G10805 (W9408, W12446);
not G10806 (W9409, W12447);
not G10807 (W9410, I822);
not G10808 (W9411, W9412);
not G10809 (W9412, W12448);
not G10810 (W9413, I823);
not G10811 (W9414, W9415);
not G10812 (W9415, W12449);
not G10813 (W9416, I306);
not G10814 (W9417, W9419);
not G10815 (W9418, W12450);
not G10816 (W9419, W12451);
not G10817 (W9420, I307);
not G10818 (W9421, W9422);
not G10819 (W9422, W12452);
not G10820 (W9423, I308);
not G10821 (W9424, W9425);
not G10822 (W9425, W12453);
nor G10823 (W9426, W12454, W12455, W12456);
not G10824 (W9427, I824);
not G10825 (W9428, W9430);
not G10826 (W9429, W12457);
not G10827 (W9430, W12458);
not G10828 (W9431, I825);
not G10829 (W9432, W9433);
not G10830 (W9433, W12459);
not G10831 (W9434, I826);
not G10832 (W9435, W9436);
not G10833 (W9436, W12460);
nor G10834 (W9437, W12461, W12462, W12463);
not G10835 (W9438, I827);
not G10836 (W9439, W9441);
not G10837 (W9440, W12464);
not G10838 (W9441, W12465);
not G10839 (W9442, I828);
not G10840 (W9443, W9444);
not G10841 (W9444, W12466);
not G10842 (W9445, I829);
not G10843 (W9446, W9447);
not G10844 (W9447, W12467);
not G10845 (W9448, I309);
not G10846 (W9449, W9451);
not G10847 (W9450, W12468);
not G10848 (W9451, W12469);
not G10849 (W9452, I310);
not G10850 (W9453, W9454);
not G10851 (W9454, W12470);
not G10852 (W9455, I311);
not G10853 (W9456, W9457);
not G10854 (W9457, W12471);
nor G10855 (W9458, W12472, W12473, W12474);
not G10856 (W9459, I830);
not G10857 (W9460, W9462);
not G10858 (W9461, W12475);
not G10859 (W9462, W12476);
not G10860 (W9463, I831);
not G10861 (W9464, W9465);
not G10862 (W9465, W12477);
not G10863 (W9466, I832);
not G10864 (W9467, W9468);
not G10865 (W9468, W12478);
not G10866 (W9469, W12479);
not G10867 (W9470, W12480);
not G10868 (W9471, W12481);
not G10869 (W9472, I805);
not G10870 (W9473, W9475);
not G10871 (W9474, I833);
not G10872 (W9475, W12482);
not G10873 (W9476, W9477);
not G10874 (W9477, W12483);
nor G10875 (W9478, W12484, W12485);
not G10876 (W9479, W9480);
not G10877 (W9480, W12486);
nor G10878 (W9481, W12487, W12488);
not G10879 (W9482, W9484);
not G10880 (W9483, I834);
not G10881 (W9484, W12489);
nor G10882 (W9485, W12490, W12491);
not G10883 (W9486, W9488);
not G10884 (W9487, I835);
not G10885 (W9488, W12492);
nor G10886 (W9489, W12493, W12494);
not G10887 (W9490, W9492);
not G10888 (W9491, I836);
not G10889 (W9492, W12495);
nor G10890 (W9493, W12496, W12497);
not G10891 (W9494, W9496);
not G10892 (W9495, I837);
not G10893 (W9496, W12498);
nor G10894 (W9497, W12499, W12500);
not G10895 (W9498, W9500);
not G10896 (W9499, I838);
not G10897 (W9500, W12501);
nor G10898 (W9501, W12502, W12503);
not G10899 (W9502, I839);
not G10900 (W9503, I840);
not G10901 (W9504, I841);
not G10902 (W9505, I842);
not G10903 (W9506, I843);
not G10904 (W9507, I844);
not G10905 (W9508, I845);
not G10906 (W9509, I846);
not G10907 (W9510, I847);
and G10908 (W9511, W12504, W12505);
not G10909 (W9512, W9514);
not G10910 (W9513, I848);
not G10911 (W9514, W12506);
not G10912 (W9515, W9517);
not G10913 (W9516, I849);
not G10914 (W9517, W12507);
not G10915 (W9518, W9520);
not G10916 (W9519, I850);
not G10917 (W9520, W12508);
not G10918 (W9521, I851);
not G10919 (W9522, W9524);
not G10920 (W9523, W12509);
not G10921 (W9524, W12510);
not G10922 (W9525, I852);
not G10923 (W9526, W9527);
not G10924 (W9527, W12511);
not G10925 (W9528, I853);
not G10926 (W9529, W9530);
not G10927 (W9530, W12512);
not G10928 (W9531, I854);
not G10929 (W9532, W9534);
not G10930 (W9533, W12513);
not G10931 (W9534, W12514);
not G10932 (W9535, I855);
not G10933 (W9536, W9537);
not G10934 (W9537, W12515);
not G10935 (W9538, I856);
not G10936 (W9539, W9540);
not G10937 (W9540, W12516);
not G10938 (W9541, I857);
not G10939 (W9542, W9544);
not G10940 (W9543, W12517);
not G10941 (W9544, W12518);
not G10942 (W9545, I858);
not G10943 (W9546, W9547);
not G10944 (W9547, W12519);
not G10945 (W9548, I859);
not G10946 (W9549, W9550);
not G10947 (W9550, W12520);
not G10948 (W9551, I860);
not G10949 (W9552, W9554);
not G10950 (W9553, W12521);
not G10951 (W9554, W12522);
not G10952 (W9555, I861);
not G10953 (W9556, W9557);
not G10954 (W9557, W12523);
not G10955 (W9558, I862);
not G10956 (W9559, W9560);
not G10957 (W9560, W12524);
not G10958 (W9561, I863);
not G10959 (W9562, W9564);
not G10960 (W9563, W12525);
not G10961 (W9564, W12526);
not G10962 (W9565, I864);
not G10963 (W9566, W9567);
not G10964 (W9567, W12527);
not G10965 (W9568, I865);
not G10966 (W9569, W9570);
not G10967 (W9570, W12528);
not G10968 (W9571, I866);
not G10969 (W9572, W9574);
not G10970 (W9573, W12529);
not G10971 (W9574, W12530);
not G10972 (W9575, I867);
not G10973 (W9576, W9577);
not G10974 (W9577, W12531);
not G10975 (W9578, I868);
not G10976 (W9579, W9580);
not G10977 (W9580, W12532);
not G10978 (W9581, I869);
not G10979 (W9582, W9584);
not G10980 (W9583, W12533);
not G10981 (W9584, W12534);
not G10982 (W9585, I870);
not G10983 (W9586, W9587);
not G10984 (W9587, W12535);
not G10985 (W9588, I871);
not G10986 (W9589, W9590);
not G10987 (W9590, W12536);
not G10988 (W9591, I872);
not G10989 (W9592, W9594);
not G10990 (W9593, W12537);
not G10991 (W9594, W12538);
not G10992 (W9595, I873);
not G10993 (W9596, W9597);
not G10994 (W9597, W12539);
not G10995 (W9598, I874);
not G10996 (W9599, W9600);
not G10997 (W9600, W12540);
not G10998 (W9601, I875);
not G10999 (W9602, W9604);
not G11000 (W9603, W12541);
not G11001 (W9604, W12542);
not G11002 (W9605, I876);
not G11003 (W9606, W9607);
not G11004 (W9607, W12543);
not G11005 (W9608, I877);
not G11006 (W9609, W9610);
not G11007 (W9610, W12544);
not G11008 (W9611, I878);
not G11009 (W9612, W9614);
not G11010 (W9613, W12545);
not G11011 (W9614, W12546);
not G11012 (W9615, I879);
not G11013 (W9616, W9617);
not G11014 (W9617, W12547);
not G11015 (W9618, I880);
not G11016 (W9619, W9620);
not G11017 (W9620, W12548);
not G11018 (W9621, I881);
not G11019 (W9622, W9624);
not G11020 (W9623, W12549);
not G11021 (W9624, W12550);
not G11022 (W9625, I882);
not G11023 (W9626, W9627);
not G11024 (W9627, W12551);
not G11025 (W9628, I883);
not G11026 (W9629, W9630);
not G11027 (W9630, W12552);
not G11028 (W9631, I884);
not G11029 (W9632, W9634);
not G11030 (W9633, W12553);
not G11031 (W9634, W12554);
not G11032 (W9635, I885);
not G11033 (W9636, W9637);
not G11034 (W9637, W12555);
not G11035 (W9638, I886);
not G11036 (W9639, W9640);
not G11037 (W9640, W12556);
not G11038 (W9641, I887);
not G11039 (W9642, W9644);
not G11040 (W9643, W12557);
not G11041 (W9644, W12558);
not G11042 (W9645, I888);
not G11043 (W9646, W9647);
not G11044 (W9647, W12559);
not G11045 (W9648, I889);
not G11046 (W9649, W9650);
not G11047 (W9650, W12560);
nor G11048 (W9651, W12561, W12562);
not G11049 (W9652, W9654);
not G11050 (W9653, I890);
not G11051 (W9654, W12563);
not G11052 (W9655, W9657);
not G11053 (W9656, I891);
not G11054 (W9657, W12564);
not G11055 (W9658, W9660);
not G11056 (W9659, I892);
not G11057 (W9660, W12565);
not G11058 (W9661, W12566);
nor G11059 (W9662, W12567, W12568);
nand G11060 (W9663, W12569, W12570);
not G11061 (W9664, W9666);
not G11062 (W9665, I329);
not G11063 (W9666, W12571);
nand G11064 (W9667, W12572, W12573, W12574);
not G11065 (W9668, W9670);
not G11066 (W9669, I326);
not G11067 (W9670, W12575);
nand G11068 (W9671, W12576, W12577);
not G11069 (W9672, W9674);
not G11070 (W9673, I323);
not G11071 (W9674, W12578);
nand G11072 (W9675, W12579, W12580);
not G11073 (W9676, W9678);
not G11074 (W9677, I320);
not G11075 (W9678, W12581);
not G11076 (W9679, W9681);
not G11077 (W9680, I330);
not G11078 (W9681, W12582);
not G11079 (W9682, W9684);
not G11080 (W9683, I331);
not G11081 (W9684, W12583);
not G11082 (W9685, W9687);
not G11083 (W9686, I327);
not G11084 (W9687, W12584);
not G11085 (W9688, W9690);
not G11086 (W9689, I328);
not G11087 (W9690, W12585);
not G11088 (W9691, W9693);
not G11089 (W9692, I324);
not G11090 (W9693, W12586);
not G11091 (W9694, W9696);
not G11092 (W9695, I325);
not G11093 (W9696, W12587);
not G11094 (W9697, W9699);
not G11095 (W9698, I321);
not G11096 (W9699, W12588);
not G11097 (W9700, W9702);
not G11098 (W9701, I322);
not G11099 (W9702, W12589);
not G11100 (W9703, I893);
not G11101 (W9704, W9706);
not G11102 (W9705, W12590);
not G11103 (W9706, W12591);
not G11104 (W9707, I894);
not G11105 (W9708, W9709);
not G11106 (W9709, W12592);
not G11107 (W9710, I895);
not G11108 (W9711, W9712);
not G11109 (W9712, W12593);
nor G11110 (W9713, W12594, W12595, W12596);
not G11111 (W9714, W9716);
not G11112 (W9715, I896);
not G11113 (W9716, W12597);
not G11114 (W9717, W9719);
not G11115 (W9718, I897);
not G11116 (W9719, W12598);
not G11117 (W9720, W9722);
not G11118 (W9721, I898);
not G11119 (W9722, W12599);
not G11120 (W9723, I899);
not G11121 (W9724, W9726);
not G11122 (W9725, W12600);
not G11123 (W9726, W12601);
not G11124 (W9727, I900);
not G11125 (W9728, W9729);
not G11126 (W9729, W12602);
not G11127 (W9730, I901);
not G11128 (W9731, W9732);
not G11129 (W9732, W12603);
not G11130 (W9733, I902);
not G11131 (W9734, W9736);
not G11132 (W9735, W12604);
not G11133 (W9736, W12605);
not G11134 (W9737, I903);
not G11135 (W9738, W9739);
not G11136 (W9739, W12606);
not G11137 (W9740, I904);
not G11138 (W9741, W9742);
not G11139 (W9742, W12607);
not G11140 (W9743, I905);
not G11141 (W9744, W9746);
not G11142 (W9745, W12608);
not G11143 (W9746, W12609);
not G11144 (W9747, I906);
not G11145 (W9748, W9749);
not G11146 (W9749, W12610);
not G11147 (W9750, I907);
not G11148 (W9751, W9752);
not G11149 (W9752, W12611);
not G11150 (W9753, W12612);
not G11151 (W9754, W9756);
not G11152 (W9755, I908);
not G11153 (W9756, W12613);
not G11154 (W9757, W9759);
not G11155 (W9758, I909);
not G11156 (W9759, W12614);
not G11157 (W9760, W9762);
not G11158 (W9761, I910);
not G11159 (W9762, W12615);
and G11160 (W9763, W12616, I902);
and G11161 (W9764, W12617, I903);
and G11162 (W9765, W12618, I904);
and G11163 (W9766, W12616, W9701);
and G11164 (W9767, W12617, W9698);
and G11165 (W9768, W12618, W9677);
and G11166 (W9769, W12616, W9695);
and G11167 (W9770, W12617, W9692);
and G11168 (W9771, W12618, W9673);
and G11169 (W9772, W12616, W9689);
and G11170 (W9773, W12617, W9686);
and G11171 (W9774, W12618, W9669);
and G11172 (W9775, W12616, W9683);
and G11173 (W9776, W12617, W9680);
and G11174 (W9777, W12618, W9665);
not G11175 (W9778, W12619);
not G11176 (W9779, W9781);
not G11177 (W9780, I911);
not G11178 (W9781, W12620);
not G11179 (W9782, W12621);
not G11180 (W9783, W9785);
not G11181 (W9784, I912);
not G11182 (W9785, W12622);
not G11183 (W9786, W12623);
not G11184 (W9787, W9789);
not G11185 (W9788, I913);
not G11186 (W9789, W12624);
not G11187 (W9790, W12625);
not G11188 (W9791, W9793);
not G11189 (W9792, I914);
not G11190 (W9793, W12626);
not G11191 (W9794, W12627);
not G11192 (W9795, W9797);
not G11193 (W9796, I915);
not G11194 (W9797, W12628);
not G11195 (W9798, W12629);
not G11196 (W9799, W9801);
not G11197 (W9800, I916);
not G11198 (W9801, W12630);
not G11199 (W9802, W12631);
not G11200 (W9803, W9805);
not G11201 (W9804, I917);
not G11202 (W9805, W12632);
not G11203 (W9806, W12633);
not G11204 (W9807, W9809);
not G11205 (W9808, I918);
not G11206 (W9809, W12634);
not G11207 (W9810, W12635);
not G11208 (W9811, W9813);
not G11209 (W9812, I919);
not G11210 (W9813, W12636);
not G11211 (W9814, W12637);
not G11212 (W9815, W9817);
not G11213 (W9816, I920);
not G11214 (W9817, W12638);
not G11215 (W9818, W9820);
not G11216 (W9819, I921);
not G11217 (W9820, W12639);
not G11218 (W9821, W9823);
not G11219 (W9822, I922);
not G11220 (W9823, W12640);
not G11221 (W9824, W9826);
not G11222 (W9825, I923);
not G11223 (W9826, W12641);
not G11224 (W9827, W9829);
not G11225 (W9828, I924);
not G11226 (W9829, W12642);
not G11227 (W9830, W9832);
not G11228 (W9831, I925);
not G11229 (W9832, W12643);
not G11230 (W9833, W9835);
not G11231 (W9834, I926);
not G11232 (W9835, W12644);
not G11233 (W9836, W9838);
not G11234 (W9837, I927);
not G11235 (W9838, W12645);
not G11236 (W9839, W9841);
not G11237 (W9840, I928);
not G11238 (W9841, W12646);
not G11239 (W9842, W9844);
not G11240 (W9843, I929);
not G11241 (W9844, W12647);
not G11242 (W9845, W9847);
not G11243 (W9846, I930);
not G11244 (W9847, W12648);
not G11245 (W9848, W9850);
not G11246 (W9849, I931);
not G11247 (W9850, W12649);
not G11248 (W9851, W9853);
not G11249 (W9852, I932);
not G11250 (W9853, W12650);
not G11251 (W9854, W9856);
not G11252 (W9855, I933);
not G11253 (W9856, W12651);
not G11254 (W9857, W9859);
not G11255 (W9858, I934);
not G11256 (W9859, W12652);
not G11257 (W9860, W9862);
not G11258 (W9861, I935);
not G11259 (W9862, W12653);
not G11260 (W9863, W9865);
not G11261 (W9864, I936);
not G11262 (W9865, W12654);
not G11263 (W9866, W9868);
not G11264 (W9867, I937);
not G11265 (W9868, W12655);
not G11266 (W9869, W9871);
not G11267 (W9870, I938);
not G11268 (W9871, W12656);
not G11269 (W9872, W9874);
not G11270 (W9873, I939);
not G11271 (W9874, W12657);
not G11272 (W9875, W9877);
not G11273 (W9876, I940);
not G11274 (W9877, W12658);
and G11275 (W9878, I941, W12659);
and G11276 (W9879, W12660, W12661);
not G11277 (W9880, W12662);
not G11278 (W9881, W12663);
not G11279 (W9882, W12664);
and G11280 (W9883, W12665, W12666);
and G11281 (W9884, I942, W12667);
and G11282 (W9885, I943, W12668);
and G11283 (W9886, W12669, W12670);
and G11284 (W9887, W12671, W12672);
and G11285 (W9888, I944, W12673);
and G11286 (W9889, I945, W12674);
and G11287 (W9890, W12675, W12676);
and G11288 (W9891, W12677, W12678);
and G11289 (W9892, I946, W12679);
and G11290 (W9893, I947, W12680);
and G11291 (W9894, W12681, W12682);
and G11292 (W9895, W12683, W12684);
and G11293 (W9896, I948, W12685);
and G11294 (W9897, I949, W12686);
and G11295 (W9898, W12687, W12688);
and G11296 (W9899, W12689, W12690);
and G11297 (W9900, I950, W12691);
and G11298 (W9901, W12692, W12693);
not G11299 (W9902, W9904);
not G11300 (W9903, I951);
not G11301 (W9904, W12694);
not G11302 (W9905, W9907);
not G11303 (W9906, I952);
not G11304 (W9907, W12695);
not G11305 (W9908, W9910);
not G11306 (W9909, I953);
not G11307 (W9910, W12696);
not G11308 (W9911, W9913);
not G11309 (W9912, I954);
not G11310 (W9913, W12697);
not G11311 (W9914, W9916);
not G11312 (W9915, I955);
not G11313 (W9916, W12698);
not G11314 (W9917, W9919);
not G11315 (W9918, I956);
not G11316 (W9919, W12699);
not G11317 (W9920, W9922);
not G11318 (W9921, I957);
not G11319 (W9922, W12700);
not G11320 (W9923, W9925);
not G11321 (W9924, I958);
not G11322 (W9925, W12701);
not G11323 (W9926, W9928);
not G11324 (W9927, I959);
not G11325 (W9928, W12702);
nand G11326 (W9929, W9786, W9798, W12703);
not G11327 (W9930, W9932);
not G11328 (W9931, I960);
not G11329 (W9932, W12704);
not G11330 (W9933, W9935);
not G11331 (W9934, I961);
not G11332 (W9935, W12705);
not G11333 (W9936, W9938);
not G11334 (W9937, I962);
not G11335 (W9938, W12706);
and G11336 (W9939, W12707, W12708);
and G11337 (W9940, W12709, W12710);
and G11338 (W9941, W12711, W12712);
and G11339 (W9942, W12713, W12714);
and G11340 (W9943, W12715, W12716);
and G11341 (W9944, W12717, W12718);
and G11342 (W9945, W12719, W12720);
and G11343 (W9946, W12721, W12722);
and G11344 (W9947, W12723, W12724);
and G11345 (W9948, W12725, W12726);
and G11346 (W9949, W12727, W12728);
and G11347 (W9950, W12729, W12730);
and G11348 (W9951, W11815, W12731);
and G11349 (W9952, W12732, W12733);
and G11350 (W9953, W12734, W12735);
and G11351 (W9954, W12736, W12737);
and G11352 (W9955, W12738, W12739);
and G11353 (W9956, W12740, W12741);
and G11354 (W9957, W12742, W12743);
not G11355 (W9958, W12744);
not G11356 (W9959, W9961);
not G11357 (W9960, I963);
not G11358 (W9961, W12745);
not G11359 (W9962, W9964);
not G11360 (W9963, I964);
not G11361 (W9964, W12746);
not G11362 (W9965, W9967);
not G11363 (W9966, I965);
not G11364 (W9967, W12747);
not G11365 (W9968, W12748);
not G11366 (W9969, W9971);
not G11367 (W9970, I966);
not G11368 (W9971, W12749);
not G11369 (W9972, W9974);
not G11370 (W9973, I967);
not G11371 (W9974, W12750);
not G11372 (W9975, W9977);
not G11373 (W9976, I968);
not G11374 (W9977, W12751);
not G11375 (W9978, W12752);
not G11376 (W9979, W9981);
not G11377 (W9980, I969);
not G11378 (W9981, W12753);
not G11379 (W9982, W9984);
not G11380 (W9983, I970);
not G11381 (W9984, W12754);
not G11382 (W9985, W9987);
not G11383 (W9986, I971);
not G11384 (W9987, W12755);
not G11385 (W9988, W12756);
not G11386 (W9989, W9991);
not G11387 (W9990, I972);
not G11388 (W9991, W12757);
not G11389 (W9992, W9994);
not G11390 (W9993, I973);
not G11391 (W9994, W12758);
not G11392 (W9995, W9997);
not G11393 (W9996, I974);
not G11394 (W9997, W12759);
not G11395 (W9998, W10000);
not G11396 (W9999, I975);
not G11397 (W10000, W12760);
not G11398 (W10001, W10003);
not G11399 (W10002, I976);
not G11400 (W10003, W12761);
not G11401 (W10004, W10006);
not G11402 (W10005, I977);
not G11403 (W10006, W12762);
not G11404 (W10007, W10009);
not G11405 (W10008, I978);
not G11406 (W10009, W12763);
not G11407 (W10010, W10012);
not G11408 (W10011, I979);
not G11409 (W10012, W12764);
not G11410 (W10013, W10015);
not G11411 (W10014, I980);
not G11412 (W10015, W12765);
not G11413 (W10016, W10018);
not G11414 (W10017, I981);
not G11415 (W10018, W12766);
not G11416 (W10019, W10021);
not G11417 (W10020, I982);
not G11418 (W10021, W12767);
not G11419 (W10022, W10024);
not G11420 (W10023, I983);
not G11421 (W10024, W12768);
not G11422 (W10025, W10027);
not G11423 (W10026, I984);
not G11424 (W10027, W12769);
not G11425 (W10028, W10030);
not G11426 (W10029, I985);
not G11427 (W10030, W12770);
not G11428 (W10031, W10033);
not G11429 (W10032, I986);
not G11430 (W10033, W12771);
not G11431 (W10034, W10036);
not G11432 (W10035, I987);
not G11433 (W10036, W12772);
not G11434 (W10037, W10039);
not G11435 (W10038, I988);
not G11436 (W10039, W12773);
not G11437 (W10040, W10042);
not G11438 (W10041, I989);
not G11439 (W10042, W12774);
not G11440 (W10043, W10045);
not G11441 (W10044, I990);
not G11442 (W10045, W12775);
not G11443 (W10046, W10048);
not G11444 (W10047, I991);
not G11445 (W10048, W12776);
not G11446 (W10049, W10051);
not G11447 (W10050, I992);
not G11448 (W10051, W12777);
not G11449 (W10052, W10054);
not G11450 (W10053, I993);
not G11451 (W10054, W12778);
not G11452 (W10055, W10057);
not G11453 (W10056, I994);
not G11454 (W10057, W12779);
not G11455 (W10058, W10060);
not G11456 (W10059, I995);
not G11457 (W10060, W12780);
not G11458 (W10061, W10063);
not G11459 (W10062, I996);
not G11460 (W10063, W12781);
not G11461 (W10064, W10066);
not G11462 (W10065, I997);
not G11463 (W10066, W12782);
not G11464 (W10067, W10069);
not G11465 (W10068, I998);
not G11466 (W10069, W12783);
not G11467 (W10070, W10072);
not G11468 (W10071, I999);
not G11469 (W10072, W12784);
not G11470 (W10073, W10075);
not G11471 (W10074, I1000);
not G11472 (W10075, W12785);
not G11473 (W10076, W10078);
not G11474 (W10077, I1001);
not G11475 (W10078, W12786);
not G11476 (W10079, W10081);
not G11477 (W10080, I1002);
not G11478 (W10081, W12787);
not G11479 (W10082, W10084);
not G11480 (W10083, I1003);
not G11481 (W10084, W12788);
not G11482 (W10085, W10087);
not G11483 (W10086, I1004);
not G11484 (W10087, W12789);
and G11485 (W10088, I332, W12790);
and G11486 (W10089, W12791, W12792);
not G11487 (W10090, W12793);
and G11488 (W10091, W12794, W12795);
and G11489 (W10092, I333, W12796);
and G11490 (W10093, I334, W12797);
and G11491 (W10094, W12798, W12799);
and G11492 (W10095, W12800, W12801);
and G11493 (W10096, I335, W12802);
and G11494 (W10097, I336, W12803);
and G11495 (W10098, W12804, W12805);
and G11496 (W10099, W12806, W12807);
and G11497 (W10100, I337, W12808);
and G11498 (W10101, I338, W12809);
and G11499 (W10102, W12810, W12811);
and G11500 (W10103, W12812, W12813);
and G11501 (W10104, I339, W12814);
and G11502 (W10105, I340, W12815);
and G11503 (W10106, W12816, W12817);
and G11504 (W10107, W12818, W12819);
and G11505 (W10108, I341, W12820);
not G11506 (W10109, I1005);
not G11507 (W10110, W10112);
not G11508 (W10111, I1006);
not G11509 (W10112, W12821);
nor G11510 (W10113, W12822, W12823);
not G11511 (W10114, W10116);
not G11512 (W10115, I1007);
not G11513 (W10116, W12824);
nor G11514 (W10117, W12825, W12826);
not G11515 (W10118, W10120);
not G11516 (W10119, I1008);
not G11517 (W10120, W12827);
nor G11518 (W10121, W12828, W12829);
not G11519 (W10122, W10124);
not G11520 (W10123, I1009);
not G11521 (W10124, W12830);
nor G11522 (W10125, W12831, W12832);
not G11523 (W10126, W10128);
not G11524 (W10127, I1010);
not G11525 (W10128, W12833);
nor G11526 (W10129, W12834, W12835);
not G11527 (W10130, W10132);
not G11528 (W10131, I1011);
not G11529 (W10132, W12836);
not G11530 (W10133, I1012);
not G11531 (W10134, W10136);
not G11532 (W10135, W12837);
not G11533 (W10136, W12838);
not G11534 (W10137, I1013);
not G11535 (W10138, W10139);
not G11536 (W10139, W12839);
not G11537 (W10140, I1014);
not G11538 (W10141, W10142);
not G11539 (W10142, W12840);
and G11540 (W10143, W10242, W8283);
and G11541 (W10144, W10243, W8280);
and G11542 (W10145, W10244, W8259);
and G11543 (W10146, W10242, W8277);
and G11544 (W10147, W10243, W8274);
and G11545 (W10148, W10244, W8255);
and G11546 (W10149, W10242, W8271);
and G11547 (W10150, W10243, W8268);
and G11548 (W10151, W10244, W8251);
and G11549 (W10152, W10242, W8265);
and G11550 (W10153, W10243, W8262);
and G11551 (W10154, W10244, W8247);
not G11552 (W10155, I1015);
not G11553 (W10156, W10158);
not G11554 (W10157, W12841);
not G11555 (W10158, W12842);
not G11556 (W10159, I1016);
not G11557 (W10160, W10161);
not G11558 (W10161, W12843);
not G11559 (W10162, I1017);
not G11560 (W10163, W10164);
not G11561 (W10164, W12844);
not G11562 (W10165, I1018);
not G11563 (W10166, W10168);
not G11564 (W10167, W12845);
not G11565 (W10168, W12846);
not G11566 (W10169, I1019);
not G11567 (W10170, W10171);
not G11568 (W10171, W12847);
not G11569 (W10172, I1020);
not G11570 (W10173, W10174);
not G11571 (W10174, W12848);
nor G11572 (W10175, W12849, W12850);
not G11573 (W10176, W10178);
not G11574 (W10177, I1021);
not G11575 (W10178, W12851);
not G11576 (W10179, I1022);
not G11577 (W10180, W10182);
not G11578 (W10181, W12852);
not G11579 (W10182, W12853);
not G11580 (W10183, I1023);
not G11581 (W10184, W10185);
not G11582 (W10185, W12854);
not G11583 (W10186, I1024);
not G11584 (W10187, W10188);
not G11585 (W10188, W12855);
not G11586 (W10189, I342);
not G11587 (W10190, W10192);
not G11588 (W10191, W12856);
not G11589 (W10192, W12857);
not G11590 (W10193, I343);
not G11591 (W10194, W10195);
not G11592 (W10195, W12858);
not G11593 (W10196, I344);
not G11594 (W10197, W10198);
not G11595 (W10198, W12859);
nor G11596 (W10199, W12860, W12861, W12862);
not G11597 (W10200, I1025);
not G11598 (W10201, W10203);
not G11599 (W10202, W12863);
not G11600 (W10203, W12864);
not G11601 (W10204, I1026);
not G11602 (W10205, W10206);
not G11603 (W10206, W12865);
not G11604 (W10207, I1027);
not G11605 (W10208, W10209);
not G11606 (W10209, W12866);
nor G11607 (W10210, W12867, W12868, W12869);
not G11608 (W10211, I1028);
not G11609 (W10212, W10214);
not G11610 (W10213, W12870);
not G11611 (W10214, W12871);
not G11612 (W10215, I1029);
not G11613 (W10216, W10217);
not G11614 (W10217, W12872);
not G11615 (W10218, I1030);
not G11616 (W10219, W10220);
not G11617 (W10220, W12873);
not G11618 (W10221, I345);
not G11619 (W10222, W10224);
not G11620 (W10223, W12874);
not G11621 (W10224, W12875);
not G11622 (W10225, I346);
not G11623 (W10226, W10227);
not G11624 (W10227, W12876);
not G11625 (W10228, I347);
not G11626 (W10229, W10230);
not G11627 (W10230, W12877);
nor G11628 (W10231, W12878, W12879, W12880);
not G11629 (W10232, I1031);
not G11630 (W10233, W10235);
not G11631 (W10234, W12881);
not G11632 (W10235, W12882);
not G11633 (W10236, I1032);
not G11634 (W10237, W10238);
not G11635 (W10238, W12883);
not G11636 (W10239, I1033);
not G11637 (W10240, W10241);
not G11638 (W10241, W12884);
not G11639 (W10242, W12885);
not G11640 (W10243, W12886);
not G11641 (W10244, W12887);
not G11642 (W10245, I1006);
not G11643 (W10246, W10248);
not G11644 (W10247, I1034);
not G11645 (W10248, W12888);
not G11646 (W10249, W10250);
not G11647 (W10250, W12889);
nor G11648 (W10251, W12890, W12891);
not G11649 (W10252, W10253);
not G11650 (W10253, W12892);
nor G11651 (W10254, W12893, W12894);
not G11652 (W10255, W10257);
not G11653 (W10256, I1035);
not G11654 (W10257, W12895);
nor G11655 (W10258, W12896, W12897);
not G11656 (W10259, W10261);
not G11657 (W10260, I1036);
not G11658 (W10261, W12898);
nor G11659 (W10262, W12899, W12900);
not G11660 (W10263, W10265);
not G11661 (W10264, I1037);
not G11662 (W10265, W12901);
nor G11663 (W10266, W12902, W12903);
not G11664 (W10267, W10269);
not G11665 (W10268, I1038);
not G11666 (W10269, W12904);
nor G11667 (W10270, W12905, W12906);
not G11668 (W10271, W10273);
not G11669 (W10272, I1039);
not G11670 (W10273, W12907);
nor G11671 (W10274, W12908, W12909);
not G11672 (W10275, I1040);
not G11673 (W10276, I1041);
not G11674 (W10277, I1042);
not G11675 (W10278, I1043);
not G11676 (W10279, I1044);
not G11677 (W10280, I1045);
not G11678 (W10281, I1046);
not G11679 (W10282, I1047);
not G11680 (W10283, I1048);
and G11681 (W10284, W12910, W12911);
not G11682 (W10285, W10287);
not G11683 (W10286, I1049);
not G11684 (W10287, W12912);
not G11685 (W10288, W10290);
not G11686 (W10289, I1050);
not G11687 (W10290, W12913);
not G11688 (W10291, W10293);
not G11689 (W10292, I1051);
not G11690 (W10293, W12914);
not G11691 (W10294, I1052);
not G11692 (W10295, W10297);
not G11693 (W10296, W12915);
not G11694 (W10297, W12916);
not G11695 (W10298, I1053);
not G11696 (W10299, W10300);
not G11697 (W10300, W12917);
not G11698 (W10301, I1054);
not G11699 (W10302, W10303);
not G11700 (W10303, W12918);
not G11701 (W10304, I1055);
not G11702 (W10305, W10307);
not G11703 (W10306, W12919);
not G11704 (W10307, W12920);
not G11705 (W10308, I1056);
not G11706 (W10309, W10310);
not G11707 (W10310, W12921);
not G11708 (W10311, I1057);
not G11709 (W10312, W10313);
not G11710 (W10313, W12922);
not G11711 (W10314, I1058);
not G11712 (W10315, W10317);
not G11713 (W10316, W12923);
not G11714 (W10317, W12924);
not G11715 (W10318, I1059);
not G11716 (W10319, W10320);
not G11717 (W10320, W12925);
not G11718 (W10321, I1060);
not G11719 (W10322, W10323);
not G11720 (W10323, W12926);
not G11721 (W10324, I1061);
not G11722 (W10325, W10327);
not G11723 (W10326, W12927);
not G11724 (W10327, W12928);
not G11725 (W10328, I1062);
not G11726 (W10329, W10330);
not G11727 (W10330, W12929);
not G11728 (W10331, I1063);
not G11729 (W10332, W10333);
not G11730 (W10333, W12930);
not G11731 (W10334, I1064);
not G11732 (W10335, W10337);
not G11733 (W10336, W12931);
not G11734 (W10337, W12932);
not G11735 (W10338, I1065);
not G11736 (W10339, W10340);
not G11737 (W10340, W12933);
not G11738 (W10341, I1066);
not G11739 (W10342, W10343);
not G11740 (W10343, W12934);
not G11741 (W10344, I1067);
not G11742 (W10345, W10347);
not G11743 (W10346, W12935);
not G11744 (W10347, W12936);
not G11745 (W10348, I1068);
not G11746 (W10349, W10350);
not G11747 (W10350, W12937);
not G11748 (W10351, I1069);
not G11749 (W10352, W10353);
not G11750 (W10353, W12938);
not G11751 (W10354, I1070);
not G11752 (W10355, W10357);
not G11753 (W10356, W12939);
not G11754 (W10357, W12940);
not G11755 (W10358, I1071);
not G11756 (W10359, W10360);
not G11757 (W10360, W12941);
not G11758 (W10361, I1072);
not G11759 (W10362, W10363);
not G11760 (W10363, W12942);
not G11761 (W10364, I1073);
not G11762 (W10365, W10367);
not G11763 (W10366, W12943);
not G11764 (W10367, W12944);
not G11765 (W10368, I1074);
not G11766 (W10369, W10370);
not G11767 (W10370, W12945);
not G11768 (W10371, I1075);
not G11769 (W10372, W10373);
not G11770 (W10373, W12946);
not G11771 (W10374, I1076);
not G11772 (W10375, W10377);
not G11773 (W10376, W12947);
not G11774 (W10377, W12948);
not G11775 (W10378, I1077);
not G11776 (W10379, W10380);
not G11777 (W10380, W12949);
not G11778 (W10381, I1078);
not G11779 (W10382, W10383);
not G11780 (W10383, W12950);
not G11781 (W10384, I1079);
not G11782 (W10385, W10387);
not G11783 (W10386, W12951);
not G11784 (W10387, W12952);
not G11785 (W10388, I1080);
not G11786 (W10389, W10390);
not G11787 (W10390, W12953);
not G11788 (W10391, I1081);
not G11789 (W10392, W10393);
not G11790 (W10393, W12954);
not G11791 (W10394, I1082);
not G11792 (W10395, W10397);
not G11793 (W10396, W12955);
not G11794 (W10397, W12956);
not G11795 (W10398, I1083);
not G11796 (W10399, W10400);
not G11797 (W10400, W12957);
not G11798 (W10401, I1084);
not G11799 (W10402, W10403);
not G11800 (W10403, W12958);
not G11801 (W10404, I1085);
not G11802 (W10405, W10407);
not G11803 (W10406, W12959);
not G11804 (W10407, W12960);
not G11805 (W10408, I1086);
not G11806 (W10409, W10410);
not G11807 (W10410, W12961);
not G11808 (W10411, I1087);
not G11809 (W10412, W10413);
not G11810 (W10413, W12962);
not G11811 (W10414, I1088);
not G11812 (W10415, W10417);
not G11813 (W10416, W12963);
not G11814 (W10417, W12964);
not G11815 (W10418, I1089);
not G11816 (W10419, W10420);
not G11817 (W10420, W12965);
not G11818 (W10421, I1090);
not G11819 (W10422, W10423);
not G11820 (W10423, W12966);
nor G11821 (W10424, W12967, W12968);
not G11822 (W10425, W10427);
not G11823 (W10426, I1091);
not G11824 (W10427, W12969);
not G11825 (W10428, W10430);
not G11826 (W10429, I1092);
not G11827 (W10430, W12970);
not G11828 (W10431, W10433);
not G11829 (W10432, I1093);
not G11830 (W10433, W12971);
not G11831 (W10434, W12972);
nor G11832 (W10435, W12973, W12974);
nand G11833 (W10436, W12975, W12976);
not G11834 (W10437, W10439);
not G11835 (W10438, I365);
not G11836 (W10439, W12977);
nand G11837 (W10440, W12978, W12979, W12980);
not G11838 (W10441, W10443);
not G11839 (W10442, I362);
not G11840 (W10443, W12981);
nand G11841 (W10444, W12982, W12983);
not G11842 (W10445, W10447);
not G11843 (W10446, I359);
not G11844 (W10447, W12984);
nand G11845 (W10448, W12985, W12986);
not G11846 (W10449, W10451);
not G11847 (W10450, I356);
not G11848 (W10451, W12987);
not G11849 (W10452, W10454);
not G11850 (W10453, I366);
not G11851 (W10454, W12988);
not G11852 (W10455, W10457);
not G11853 (W10456, I367);
not G11854 (W10457, W12989);
not G11855 (W10458, W10460);
not G11856 (W10459, I363);
not G11857 (W10460, W12990);
not G11858 (W10461, W10463);
not G11859 (W10462, I364);
not G11860 (W10463, W12991);
not G11861 (W10464, W10466);
not G11862 (W10465, I360);
not G11863 (W10466, W12992);
not G11864 (W10467, W10469);
not G11865 (W10468, I361);
not G11866 (W10469, W12993);
not G11867 (W10470, W10472);
not G11868 (W10471, I357);
not G11869 (W10472, W12994);
not G11870 (W10473, W10475);
not G11871 (W10474, I358);
not G11872 (W10475, W12995);
not G11873 (W10476, I1094);
not G11874 (W10477, W10479);
not G11875 (W10478, W12996);
not G11876 (W10479, W12997);
not G11877 (W10480, I1095);
not G11878 (W10481, W10482);
not G11879 (W10482, W12998);
not G11880 (W10483, I1096);
not G11881 (W10484, W10485);
not G11882 (W10485, W12999);
nor G11883 (W10486, W13000, W13001, W13002);
not G11884 (W10487, W10489);
not G11885 (W10488, I1097);
not G11886 (W10489, W13003);
not G11887 (W10490, W10492);
not G11888 (W10491, I1098);
not G11889 (W10492, W13004);
not G11890 (W10493, W10495);
not G11891 (W10494, I1099);
not G11892 (W10495, W13005);
not G11893 (W10496, I1100);
not G11894 (W10497, W10499);
not G11895 (W10498, W13006);
not G11896 (W10499, W13007);
not G11897 (W10500, I1101);
not G11898 (W10501, W10502);
not G11899 (W10502, W13008);
not G11900 (W10503, I1102);
not G11901 (W10504, W10505);
not G11902 (W10505, W13009);
not G11903 (W10506, I1103);
not G11904 (W10507, W10509);
not G11905 (W10508, W13010);
not G11906 (W10509, W13011);
not G11907 (W10510, I1104);
not G11908 (W10511, W10512);
not G11909 (W10512, W13012);
not G11910 (W10513, I1105);
not G11911 (W10514, W10515);
not G11912 (W10515, W13013);
not G11913 (W10516, I1106);
not G11914 (W10517, W10519);
not G11915 (W10518, W13014);
not G11916 (W10519, W13015);
not G11917 (W10520, I1107);
not G11918 (W10521, W10522);
not G11919 (W10522, W13016);
not G11920 (W10523, I1108);
not G11921 (W10524, W10525);
not G11922 (W10525, W13017);
not G11923 (W10526, W13018);
not G11924 (W10527, W10529);
not G11925 (W10528, I1109);
not G11926 (W10529, W13019);
not G11927 (W10530, W10532);
not G11928 (W10531, I1110);
not G11929 (W10532, W13020);
not G11930 (W10533, W10535);
not G11931 (W10534, I1111);
not G11932 (W10535, W13021);
and G11933 (W10536, W13022, I1103);
and G11934 (W10537, W13023, I1104);
and G11935 (W10538, W13024, I1105);
and G11936 (W10539, W13022, W10474);
and G11937 (W10540, W13023, W10471);
and G11938 (W10541, W13024, W10450);
and G11939 (W10542, W13022, W10468);
and G11940 (W10543, W13023, W10465);
and G11941 (W10544, W13024, W10446);
and G11942 (W10545, W13022, W10462);
and G11943 (W10546, W13023, W10459);
and G11944 (W10547, W13024, W10442);
and G11945 (W10548, W13022, W10456);
and G11946 (W10549, W13023, W10453);
and G11947 (W10550, W13024, W10438);
not G11948 (W10551, W13025);
not G11949 (W10552, W10554);
not G11950 (W10553, I1112);
not G11951 (W10554, W13026);
not G11952 (W10555, W13027);
not G11953 (W10556, W10558);
not G11954 (W10557, I1113);
not G11955 (W10558, W13028);
not G11956 (W10559, W13029);
not G11957 (W10560, W10562);
not G11958 (W10561, I1114);
not G11959 (W10562, W13030);
not G11960 (W10563, W13031);
not G11961 (W10564, W10566);
not G11962 (W10565, I1115);
not G11963 (W10566, W13032);
not G11964 (W10567, W13033);
not G11965 (W10568, W10570);
not G11966 (W10569, I1116);
not G11967 (W10570, W13034);
not G11968 (W10571, W13035);
not G11969 (W10572, W10574);
not G11970 (W10573, I1117);
not G11971 (W10574, W13036);
not G11972 (W10575, W13037);
not G11973 (W10576, W10578);
not G11974 (W10577, I1118);
not G11975 (W10578, W13038);
not G11976 (W10579, W13039);
not G11977 (W10580, W10582);
not G11978 (W10581, I1119);
not G11979 (W10582, W13040);
not G11980 (W10583, W13041);
not G11981 (W10584, W10586);
not G11982 (W10585, I1120);
not G11983 (W10586, W13042);
not G11984 (W10587, W13043);
not G11985 (W10588, W10590);
not G11986 (W10589, I1121);
not G11987 (W10590, W13044);
not G11988 (W10591, W10593);
not G11989 (W10592, I1122);
not G11990 (W10593, W13045);
not G11991 (W10594, W10596);
not G11992 (W10595, I1123);
not G11993 (W10596, W13046);
not G11994 (W10597, W10599);
not G11995 (W10598, I1124);
not G11996 (W10599, W13047);
not G11997 (W10600, W10602);
not G11998 (W10601, I1125);
not G11999 (W10602, W13048);
not G12000 (W10603, W10605);
not G12001 (W10604, I1126);
not G12002 (W10605, W13049);
not G12003 (W10606, W10608);
not G12004 (W10607, I1127);
not G12005 (W10608, W13050);
not G12006 (W10609, W10611);
not G12007 (W10610, I1128);
not G12008 (W10611, W13051);
not G12009 (W10612, W10614);
not G12010 (W10613, I1129);
not G12011 (W10614, W13052);
not G12012 (W10615, W10617);
not G12013 (W10616, I1130);
not G12014 (W10617, W13053);
not G12015 (W10618, W10620);
not G12016 (W10619, I1131);
not G12017 (W10620, W13054);
not G12018 (W10621, W10623);
not G12019 (W10622, I1132);
not G12020 (W10623, W13055);
not G12021 (W10624, W10626);
not G12022 (W10625, I1133);
not G12023 (W10626, W13056);
not G12024 (W10627, W10629);
not G12025 (W10628, I1134);
not G12026 (W10629, W13057);
not G12027 (W10630, W10632);
not G12028 (W10631, I1135);
not G12029 (W10632, W13058);
not G12030 (W10633, W10635);
not G12031 (W10634, I1136);
not G12032 (W10635, W13059);
not G12033 (W10636, W10638);
not G12034 (W10637, I1137);
not G12035 (W10638, W13060);
not G12036 (W10639, W10641);
not G12037 (W10640, I1138);
not G12038 (W10641, W13061);
not G12039 (W10642, W10644);
not G12040 (W10643, I1139);
not G12041 (W10644, W13062);
not G12042 (W10645, W10647);
not G12043 (W10646, I1140);
not G12044 (W10647, W13063);
not G12045 (W10648, W10650);
not G12046 (W10649, I1141);
not G12047 (W10650, W13064);
and G12048 (W10651, I1142, W13065);
and G12049 (W10652, W13066, W13067);
not G12050 (W10653, W13068);
not G12051 (W10654, W13069);
not G12052 (W10655, W13070);
and G12053 (W10656, W13071, W13072);
and G12054 (W10657, I1143, W13073);
and G12055 (W10658, I1144, W13074);
and G12056 (W10659, W13075, W13076);
and G12057 (W10660, W13077, W13078);
and G12058 (W10661, I1145, W13079);
and G12059 (W10662, I1146, W13080);
and G12060 (W10663, W13081, W13082);
and G12061 (W10664, W13083, W13084);
and G12062 (W10665, I1147, W13085);
and G12063 (W10666, I1148, W13086);
and G12064 (W10667, W13087, W13088);
and G12065 (W10668, W13089, W13090);
and G12066 (W10669, I1149, W13091);
and G12067 (W10670, I1150, W13092);
and G12068 (W10671, W13093, W13094);
and G12069 (W10672, W13095, W13096);
and G12070 (W10673, I1151, W13097);
and G12071 (W10674, W13098, W13099);
not G12072 (W10675, W10677);
not G12073 (W10676, I1152);
not G12074 (W10677, W13100);
not G12075 (W10678, W10680);
not G12076 (W10679, I1153);
not G12077 (W10680, W13101);
not G12078 (W10681, W10683);
not G12079 (W10682, I1154);
not G12080 (W10683, W13102);
not G12081 (W10684, W10686);
not G12082 (W10685, I1155);
not G12083 (W10686, W13103);
not G12084 (W10687, W10689);
not G12085 (W10688, I1156);
not G12086 (W10689, W13104);
not G12087 (W10690, W10692);
not G12088 (W10691, I1157);
not G12089 (W10692, W13105);
not G12090 (W10693, W10695);
not G12091 (W10694, I1158);
not G12092 (W10695, W13106);
not G12093 (W10696, W10698);
not G12094 (W10697, I1159);
not G12095 (W10698, W13107);
not G12096 (W10699, W10701);
not G12097 (W10700, I1160);
not G12098 (W10701, W13108);
nand G12099 (W10702, W10555, W10567, W13109);
not G12100 (W10703, W10705);
not G12101 (W10704, I1161);
not G12102 (W10705, W13110);
not G12103 (W10706, W10708);
not G12104 (W10707, I1162);
not G12105 (W10708, W13111);
not G12106 (W10709, W10711);
not G12107 (W10710, I1163);
not G12108 (W10711, W13112);
and G12109 (W10712, W13113, W13114);
and G12110 (W10713, W13115, W13116);
and G12111 (W10714, W13117, W13118);
and G12112 (W10715, W13119, W13120);
and G12113 (W10716, W13121, W13122);
and G12114 (W10717, W13123, W13124);
and G12115 (W10718, W13125, W13126);
and G12116 (W10719, W13127, W13128);
and G12117 (W10720, W13129, W13130);
and G12118 (W10721, W13131, W13132);
and G12119 (W10722, W13133, W13134);
and G12120 (W10723, W13135, W13136);
and G12121 (W10724, W11788, W13137);
and G12122 (W10725, W13138, W13139);
and G12123 (W10726, W13140, W13141);
and G12124 (W10727, W13142, W13143);
and G12125 (W10728, W13144, W13145);
and G12126 (W10729, W13146, W13147);
and G12127 (W10730, W13148, W13149);
not G12128 (W10731, W13150);
not G12129 (W10732, W10734);
not G12130 (W10733, I1164);
not G12131 (W10734, W13151);
not G12132 (W10735, W10737);
not G12133 (W10736, I1165);
not G12134 (W10737, W13152);
not G12135 (W10738, W10740);
not G12136 (W10739, I1166);
not G12137 (W10740, W13153);
not G12138 (W10741, W13154);
not G12139 (W10742, W10744);
not G12140 (W10743, I1167);
not G12141 (W10744, W13155);
not G12142 (W10745, W10747);
not G12143 (W10746, I1168);
not G12144 (W10747, W13156);
not G12145 (W10748, W10750);
not G12146 (W10749, I1169);
not G12147 (W10750, W13157);
not G12148 (W10751, W13158);
not G12149 (W10752, W10754);
not G12150 (W10753, I1170);
not G12151 (W10754, W13159);
not G12152 (W10755, W10757);
not G12153 (W10756, I1171);
not G12154 (W10757, W13160);
not G12155 (W10758, W10760);
not G12156 (W10759, I1172);
not G12157 (W10760, W13161);
not G12158 (W10761, W13162);
not G12159 (W10762, W10764);
not G12160 (W10763, I1173);
not G12161 (W10764, W13163);
not G12162 (W10765, W10767);
not G12163 (W10766, I1174);
not G12164 (W10767, W13164);
not G12165 (W10768, W10770);
not G12166 (W10769, I1175);
not G12167 (W10770, W13165);
not G12168 (W10771, W10773);
not G12169 (W10772, I1176);
not G12170 (W10773, W13166);
not G12171 (W10774, W10776);
not G12172 (W10775, I1177);
not G12173 (W10776, W13167);
not G12174 (W10777, W10779);
not G12175 (W10778, I1178);
not G12176 (W10779, W13168);
not G12177 (W10780, W10782);
not G12178 (W10781, I1179);
not G12179 (W10782, W13169);
not G12180 (W10783, W10785);
not G12181 (W10784, I1180);
not G12182 (W10785, W13170);
not G12183 (W10786, W10788);
not G12184 (W10787, I1181);
not G12185 (W10788, W13171);
not G12186 (W10789, W10791);
not G12187 (W10790, I1182);
not G12188 (W10791, W13172);
not G12189 (W10792, W10794);
not G12190 (W10793, I1183);
not G12191 (W10794, W13173);
not G12192 (W10795, W10797);
not G12193 (W10796, I1184);
not G12194 (W10797, W13174);
not G12195 (W10798, W10800);
not G12196 (W10799, I1185);
not G12197 (W10800, W13175);
not G12198 (W10801, W10803);
not G12199 (W10802, I1186);
not G12200 (W10803, W13176);
not G12201 (W10804, W10806);
not G12202 (W10805, I1187);
not G12203 (W10806, W13177);
not G12204 (W10807, W10809);
not G12205 (W10808, I1188);
not G12206 (W10809, W13178);
not G12207 (W10810, W10812);
not G12208 (W10811, I1189);
not G12209 (W10812, W13179);
not G12210 (W10813, W10815);
not G12211 (W10814, I1190);
not G12212 (W10815, W13180);
not G12213 (W10816, W10818);
not G12214 (W10817, I1191);
not G12215 (W10818, W13181);
not G12216 (W10819, W10821);
not G12217 (W10820, I1192);
not G12218 (W10821, W13182);
not G12219 (W10822, W10824);
not G12220 (W10823, I1193);
not G12221 (W10824, W13183);
not G12222 (W10825, W10827);
not G12223 (W10826, I1194);
not G12224 (W10827, W13184);
not G12225 (W10828, W10830);
not G12226 (W10829, I1195);
not G12227 (W10830, W13185);
not G12228 (W10831, W10833);
not G12229 (W10832, I1196);
not G12230 (W10833, W13186);
not G12231 (W10834, W10836);
not G12232 (W10835, I1197);
not G12233 (W10836, W13187);
not G12234 (W10837, W10839);
not G12235 (W10838, I1198);
not G12236 (W10839, W13188);
not G12237 (W10840, W10842);
not G12238 (W10841, I1199);
not G12239 (W10842, W13189);
not G12240 (W10843, W10845);
not G12241 (W10844, I1200);
not G12242 (W10845, W13190);
not G12243 (W10846, W10848);
not G12244 (W10847, I1201);
not G12245 (W10848, W13191);
not G12246 (W10849, W10851);
not G12247 (W10850, I1202);
not G12248 (W10851, W13192);
not G12249 (W10852, W10854);
not G12250 (W10853, I1203);
not G12251 (W10854, W13193);
not G12252 (W10855, W10857);
not G12253 (W10856, I1204);
not G12254 (W10857, W13194);
not G12255 (W10858, W10860);
not G12256 (W10859, I1205);
not G12257 (W10860, W13195);
and G12258 (W10861, I368, W13196);
and G12259 (W10862, W13197, W13198);
not G12260 (W10863, W13199);
and G12261 (W10864, W13200, W13201);
and G12262 (W10865, I369, W13202);
and G12263 (W10866, I370, W13203);
and G12264 (W10867, W13204, W13205);
and G12265 (W10868, W13206, W13207);
and G12266 (W10869, I371, W13208);
and G12267 (W10870, I372, W13209);
and G12268 (W10871, W13210, W13211);
and G12269 (W10872, W13212, W13213);
and G12270 (W10873, I373, W13214);
and G12271 (W10874, I374, W13215);
and G12272 (W10875, W13216, W13217);
and G12273 (W10876, W13218, W13219);
and G12274 (W10877, I375, W13220);
and G12275 (W10878, I376, W13221);
and G12276 (W10879, W13222, W13223);
and G12277 (W10880, W13224, W13225);
and G12278 (W10881, I377, W13226);
not G12279 (W10882, I1206);
not G12280 (W10883, W10885);
not G12281 (W10884, I1207);
not G12282 (W10885, W13227);
nor G12283 (W10886, W13228, W13229);
not G12284 (W10887, W10889);
not G12285 (W10888, I1208);
not G12286 (W10889, W13230);
not G12287 (W10890, W13231);
not G12288 (W10891, W10893);
not G12289 (W10892, I1209);
not G12290 (W10893, W13232);
not G12291 (W10894, W13233);
not G12292 (W10895, W10897);
not G12293 (W10896, I1210);
not G12294 (W10897, W13234);
not G12295 (W10898, W13235);
not G12296 (W10899, W10901);
not G12297 (W10900, I1211);
not G12298 (W10901, W13236);
not G12299 (W10902, W13237);
not G12300 (W10903, W10905);
not G12301 (W10904, I1212);
not G12302 (W10905, W13238);
not G12303 (W10906, I1213);
not G12304 (W10907, W10909);
not G12305 (W10908, W13239);
not G12306 (W10909, W13240);
not G12307 (W10910, I1214);
not G12308 (W10911, W10912);
not G12309 (W10912, W13241);
not G12310 (W10913, I1215);
not G12311 (W10914, W10915);
not G12312 (W10915, W13242);
and G12313 (W10916, W11015, W8239);
and G12314 (W10917, W11016, W8236);
and G12315 (W10918, W11017, W8215);
and G12316 (W10919, W11015, W8233);
and G12317 (W10920, W11016, W8230);
and G12318 (W10921, W11017, W8211);
and G12319 (W10922, W11015, W8227);
and G12320 (W10923, W11016, W8224);
and G12321 (W10924, W11017, W8207);
and G12322 (W10925, W11015, W8221);
and G12323 (W10926, W11016, W8218);
and G12324 (W10927, W11017, W8203);
not G12325 (W10928, I1216);
not G12326 (W10929, W10931);
not G12327 (W10930, W13243);
not G12328 (W10931, W13244);
not G12329 (W10932, I1217);
not G12330 (W10933, W10934);
not G12331 (W10934, W13245);
not G12332 (W10935, I1218);
not G12333 (W10936, W10937);
not G12334 (W10937, W13246);
not G12335 (W10938, I1219);
not G12336 (W10939, W10941);
not G12337 (W10940, W13247);
not G12338 (W10941, W13248);
not G12339 (W10942, I1220);
not G12340 (W10943, W10944);
not G12341 (W10944, W13249);
not G12342 (W10945, I1221);
not G12343 (W10946, W10947);
not G12344 (W10947, W13250);
not G12345 (W10948, W13251);
not G12346 (W10949, W10951);
not G12347 (W10950, I1222);
not G12348 (W10951, W13252);
not G12349 (W10952, I1223);
not G12350 (W10953, W10955);
not G12351 (W10954, W13253);
not G12352 (W10955, W13254);
not G12353 (W10956, I1224);
not G12354 (W10957, W10958);
not G12355 (W10958, W13255);
not G12356 (W10959, I1225);
not G12357 (W10960, W10961);
not G12358 (W10961, W13256);
not G12359 (W10962, I378);
not G12360 (W10963, W10965);
not G12361 (W10964, W13257);
not G12362 (W10965, W13258);
not G12363 (W10966, I379);
not G12364 (W10967, W10968);
not G12365 (W10968, W13259);
not G12366 (W10969, I380);
not G12367 (W10970, W10971);
not G12368 (W10971, W13260);
nor G12369 (W10972, W13261, W13262, W13263);
not G12370 (W10973, I1226);
not G12371 (W10974, W10976);
not G12372 (W10975, W13264);
not G12373 (W10976, W13265);
not G12374 (W10977, I1227);
not G12375 (W10978, W10979);
not G12376 (W10979, W13266);
not G12377 (W10980, I1228);
not G12378 (W10981, W10982);
not G12379 (W10982, W13267);
nor G12380 (W10983, W13268, W13269, W13270);
not G12381 (W10984, I1229);
not G12382 (W10985, W10987);
not G12383 (W10986, W13271);
not G12384 (W10987, W13272);
not G12385 (W10988, I1230);
not G12386 (W10989, W10990);
not G12387 (W10990, W13273);
not G12388 (W10991, I1231);
not G12389 (W10992, W10993);
not G12390 (W10993, W13274);
not G12391 (W10994, I381);
not G12392 (W10995, W10997);
not G12393 (W10996, W13275);
not G12394 (W10997, W13276);
not G12395 (W10998, I382);
not G12396 (W10999, W11000);
not G12397 (W11000, W13277);
not G12398 (W11001, I383);
not G12399 (W11002, W11003);
not G12400 (W11003, W13278);
nor G12401 (W11004, W13279, W13280, W13281);
not G12402 (W11005, I1232);
not G12403 (W11006, W11008);
not G12404 (W11007, W13282);
not G12405 (W11008, W13283);
not G12406 (W11009, I1233);
not G12407 (W11010, W11011);
not G12408 (W11011, W13284);
not G12409 (W11012, I1234);
not G12410 (W11013, W11014);
not G12411 (W11014, W13285);
not G12412 (W11015, W13286);
not G12413 (W11016, W13287);
not G12414 (W11017, W13288);
not G12415 (W11018, I1207);
not G12416 (W11019, W11021);
not G12417 (W11020, I1235);
not G12418 (W11021, W13289);
not G12419 (W11022, W11023);
not G12420 (W11023, W13290);
not G12421 (W11024, W13291);
not G12422 (W11025, W11026);
not G12423 (W11026, W13292);
not G12424 (W11027, W13293);
not G12425 (W11028, W11030);
not G12426 (W11029, I1236);
not G12427 (W11030, W13294);
not G12428 (W11031, W13295);
not G12429 (W11032, W11034);
not G12430 (W11033, I1237);
not G12431 (W11034, W13296);
not G12432 (W11035, W13297);
not G12433 (W11036, W11038);
not G12434 (W11037, I1238);
not G12435 (W11038, W13298);
not G12436 (W11039, W13299);
not G12437 (W11040, W11042);
not G12438 (W11041, I1239);
not G12439 (W11042, W13300);
not G12440 (W11043, W13301);
not G12441 (W11044, W11046);
not G12442 (W11045, I1240);
not G12443 (W11046, W13302);
nor G12444 (W11047, W13303, W13304);
not G12445 (W11048, I1241);
not G12446 (W11049, I1242);
not G12447 (W11050, I1243);
not G12448 (W11051, I1244);
not G12449 (W11052, I1245);
not G12450 (W11053, I1246);
not G12451 (W11054, I1247);
not G12452 (W11055, I1248);
not G12453 (W11056, I1249);
and G12454 (W11057, W13305, W13306);
not G12455 (W11058, W11060);
not G12456 (W11059, I1250);
not G12457 (W11060, W13307);
not G12458 (W11061, W11063);
not G12459 (W11062, I1251);
not G12460 (W11063, W13308);
not G12461 (W11064, W11066);
not G12462 (W11065, I1252);
not G12463 (W11066, W13309);
not G12464 (W11067, I1253);
not G12465 (W11068, W11070);
not G12466 (W11069, W13310);
not G12467 (W11070, W13311);
not G12468 (W11071, I1254);
not G12469 (W11072, W11073);
not G12470 (W11073, W13312);
not G12471 (W11074, I1255);
not G12472 (W11075, W11076);
not G12473 (W11076, W13313);
not G12474 (W11077, I1256);
not G12475 (W11078, W11080);
not G12476 (W11079, W13314);
not G12477 (W11080, W13315);
not G12478 (W11081, I1257);
not G12479 (W11082, W11083);
not G12480 (W11083, W13316);
not G12481 (W11084, I1258);
not G12482 (W11085, W11086);
not G12483 (W11086, W13317);
not G12484 (W11087, I1259);
not G12485 (W11088, W11090);
not G12486 (W11089, W13318);
not G12487 (W11090, W13319);
not G12488 (W11091, I1260);
not G12489 (W11092, W11093);
not G12490 (W11093, W13320);
not G12491 (W11094, I1261);
not G12492 (W11095, W11096);
not G12493 (W11096, W13321);
not G12494 (W11097, I1262);
not G12495 (W11098, W11100);
not G12496 (W11099, W13322);
not G12497 (W11100, W13323);
not G12498 (W11101, I1263);
not G12499 (W11102, W11103);
not G12500 (W11103, W13324);
not G12501 (W11104, I1264);
not G12502 (W11105, W11106);
not G12503 (W11106, W13325);
not G12504 (W11107, I1265);
not G12505 (W11108, W11110);
not G12506 (W11109, W13326);
not G12507 (W11110, W13327);
not G12508 (W11111, I1266);
not G12509 (W11112, W11113);
not G12510 (W11113, W13328);
not G12511 (W11114, I1267);
not G12512 (W11115, W11116);
not G12513 (W11116, W13329);
not G12514 (W11117, I1268);
not G12515 (W11118, W11120);
not G12516 (W11119, W13330);
not G12517 (W11120, W13331);
not G12518 (W11121, I1269);
not G12519 (W11122, W11123);
not G12520 (W11123, W13332);
not G12521 (W11124, I1270);
not G12522 (W11125, W11126);
not G12523 (W11126, W13333);
not G12524 (W11127, I1271);
not G12525 (W11128, W11130);
not G12526 (W11129, W13334);
not G12527 (W11130, W13335);
not G12528 (W11131, I1272);
not G12529 (W11132, W11133);
not G12530 (W11133, W13336);
not G12531 (W11134, I1273);
not G12532 (W11135, W11136);
not G12533 (W11136, W13337);
not G12534 (W11137, I1274);
not G12535 (W11138, W11140);
not G12536 (W11139, W13338);
not G12537 (W11140, W13339);
not G12538 (W11141, I1275);
not G12539 (W11142, W11143);
not G12540 (W11143, W13340);
not G12541 (W11144, I1276);
not G12542 (W11145, W11146);
not G12543 (W11146, W13341);
not G12544 (W11147, I1277);
not G12545 (W11148, W11150);
not G12546 (W11149, W13342);
not G12547 (W11150, W13343);
not G12548 (W11151, I1278);
not G12549 (W11152, W11153);
not G12550 (W11153, W13344);
not G12551 (W11154, I1279);
not G12552 (W11155, W11156);
not G12553 (W11156, W13345);
not G12554 (W11157, I1280);
not G12555 (W11158, W11160);
not G12556 (W11159, W13346);
not G12557 (W11160, W13347);
not G12558 (W11161, I1281);
not G12559 (W11162, W11163);
not G12560 (W11163, W13348);
not G12561 (W11164, I1282);
not G12562 (W11165, W11166);
not G12563 (W11166, W13349);
not G12564 (W11167, I1283);
not G12565 (W11168, W11170);
not G12566 (W11169, W13350);
not G12567 (W11170, W13351);
not G12568 (W11171, I1284);
not G12569 (W11172, W11173);
not G12570 (W11173, W13352);
not G12571 (W11174, I1285);
not G12572 (W11175, W11176);
not G12573 (W11176, W13353);
not G12574 (W11177, I1286);
not G12575 (W11178, W11180);
not G12576 (W11179, W13354);
not G12577 (W11180, W13355);
not G12578 (W11181, I1287);
not G12579 (W11182, W11183);
not G12580 (W11183, W13356);
not G12581 (W11184, I1288);
not G12582 (W11185, W11186);
not G12583 (W11186, W13357);
not G12584 (W11187, I1289);
not G12585 (W11188, W11190);
not G12586 (W11189, W13358);
not G12587 (W11190, W13359);
not G12588 (W11191, I1290);
not G12589 (W11192, W11193);
not G12590 (W11193, W13360);
not G12591 (W11194, I1291);
not G12592 (W11195, W11196);
not G12593 (W11196, W13361);
nor G12594 (W11197, W13362, W13363);
not G12595 (W11198, W11200);
not G12596 (W11199, I1292);
not G12597 (W11200, W13364);
not G12598 (W11201, W11203);
not G12599 (W11202, I1293);
not G12600 (W11203, W13365);
not G12601 (W11204, W11206);
not G12602 (W11205, I1294);
not G12603 (W11206, W13366);
not G12604 (W11207, W13367);
nor G12605 (W11208, W13368, W13369);
nand G12606 (W11209, W13370, W13371);
not G12607 (W11210, W11212);
not G12608 (W11211, I401);
not G12609 (W11212, W13372);
nand G12610 (W11213, W13373, W13374, W13375);
not G12611 (W11214, W11216);
not G12612 (W11215, I398);
not G12613 (W11216, W13376);
nand G12614 (W11217, W13377, W13378);
not G12615 (W11218, W11220);
not G12616 (W11219, I395);
not G12617 (W11220, W13379);
nand G12618 (W11221, W13380, W13381);
not G12619 (W11222, W11224);
not G12620 (W11223, I392);
not G12621 (W11224, W13382);
not G12622 (W11225, W11227);
not G12623 (W11226, I402);
not G12624 (W11227, W13383);
not G12625 (W11228, W11230);
not G12626 (W11229, I403);
not G12627 (W11230, W13384);
not G12628 (W11231, W11233);
not G12629 (W11232, I399);
not G12630 (W11233, W13385);
not G12631 (W11234, W11236);
not G12632 (W11235, I400);
not G12633 (W11236, W13386);
not G12634 (W11237, W11239);
not G12635 (W11238, I396);
not G12636 (W11239, W13387);
not G12637 (W11240, W11242);
not G12638 (W11241, I397);
not G12639 (W11242, W13388);
not G12640 (W11243, W11245);
not G12641 (W11244, I393);
not G12642 (W11245, W13389);
not G12643 (W11246, W11248);
not G12644 (W11247, I394);
not G12645 (W11248, W13390);
not G12646 (W11249, I1295);
not G12647 (W11250, W11252);
not G12648 (W11251, W13391);
not G12649 (W11252, W13392);
not G12650 (W11253, I1296);
not G12651 (W11254, W11255);
not G12652 (W11255, W13393);
not G12653 (W11256, I1297);
not G12654 (W11257, W11258);
not G12655 (W11258, W13394);
nor G12656 (W11259, W13395, W13396, W13397);
not G12657 (W11260, W11262);
not G12658 (W11261, I1298);
not G12659 (W11262, W13398);
not G12660 (W11263, W11265);
not G12661 (W11264, I1299);
not G12662 (W11265, W13399);
not G12663 (W11266, W11268);
not G12664 (W11267, I1300);
not G12665 (W11268, W13400);
not G12666 (W11269, I1301);
not G12667 (W11270, W11272);
not G12668 (W11271, W13401);
not G12669 (W11272, W13402);
not G12670 (W11273, I1302);
not G12671 (W11274, W11275);
not G12672 (W11275, W13403);
not G12673 (W11276, I1303);
not G12674 (W11277, W11278);
not G12675 (W11278, W13404);
not G12676 (W11279, I1304);
not G12677 (W11280, W11282);
not G12678 (W11281, W13405);
not G12679 (W11282, W13406);
not G12680 (W11283, I1305);
not G12681 (W11284, W11285);
not G12682 (W11285, W13407);
not G12683 (W11286, I1306);
not G12684 (W11287, W11288);
not G12685 (W11288, W13408);
not G12686 (W11289, I1307);
not G12687 (W11290, W11292);
not G12688 (W11291, W13409);
not G12689 (W11292, W13410);
not G12690 (W11293, I1308);
not G12691 (W11294, W11295);
not G12692 (W11295, W13411);
not G12693 (W11296, I1309);
not G12694 (W11297, W11298);
not G12695 (W11298, W13412);
not G12696 (W11299, W13413);
not G12697 (W11300, W11302);
not G12698 (W11301, I1310);
not G12699 (W11302, W13414);
not G12700 (W11303, W11305);
not G12701 (W11304, I1311);
not G12702 (W11305, W13415);
not G12703 (W11306, W11308);
not G12704 (W11307, I1312);
not G12705 (W11308, W13416);
and G12706 (W11309, W13417, I1304);
and G12707 (W11310, W13418, I1305);
and G12708 (W11311, W13419, I1306);
and G12709 (W11312, W13417, W11247);
and G12710 (W11313, W13418, W11244);
and G12711 (W11314, W13419, W11223);
and G12712 (W11315, W13417, W11241);
and G12713 (W11316, W13418, W11238);
and G12714 (W11317, W13419, W11219);
and G12715 (W11318, W13417, W11235);
and G12716 (W11319, W13418, W11232);
and G12717 (W11320, W13419, W11215);
and G12718 (W11321, W13417, W11229);
and G12719 (W11322, W13418, W11226);
and G12720 (W11323, W13419, W11211);
not G12721 (W11324, W13420);
not G12722 (W11325, W11327);
not G12723 (W11326, I1313);
not G12724 (W11327, W13421);
not G12725 (W11328, W13422);
not G12726 (W11329, W11331);
not G12727 (W11330, I1314);
not G12728 (W11331, W13423);
not G12729 (W11332, W13424);
not G12730 (W11333, W11335);
not G12731 (W11334, I1315);
not G12732 (W11335, W13425);
not G12733 (W11336, W13426);
not G12734 (W11337, W11339);
not G12735 (W11338, I1316);
not G12736 (W11339, W13427);
not G12737 (W11340, W13428);
not G12738 (W11341, W11343);
not G12739 (W11342, I1317);
not G12740 (W11343, W13429);
not G12741 (W11344, W13430);
not G12742 (W11345, W11347);
not G12743 (W11346, I1318);
not G12744 (W11347, W13431);
not G12745 (W11348, W13432);
not G12746 (W11349, W11351);
not G12747 (W11350, I1319);
not G12748 (W11351, W13433);
not G12749 (W11352, W13434);
not G12750 (W11353, W11355);
not G12751 (W11354, I1320);
not G12752 (W11355, W13435);
not G12753 (W11356, W13436);
not G12754 (W11357, W11359);
not G12755 (W11358, I1321);
not G12756 (W11359, W13437);
not G12757 (W11360, W11362);
not G12758 (W11361, I1322);
not G12759 (W11362, W13438);
not G12760 (W11363, W13439);
not G12761 (W11364, W11366);
not G12762 (W11365, I1323);
not G12763 (W11366, W13440);
not G12764 (W11367, W11369);
not G12765 (W11368, I1324);
not G12766 (W11369, W13441);
not G12767 (W11370, W11372);
not G12768 (W11371, I1325);
not G12769 (W11372, W13442);
not G12770 (W11373, W11375);
not G12771 (W11374, I1326);
not G12772 (W11375, W13443);
not G12773 (W11376, W11378);
not G12774 (W11377, I1327);
not G12775 (W11378, W13444);
not G12776 (W11379, W11381);
not G12777 (W11380, I1328);
not G12778 (W11381, W13445);
not G12779 (W11382, W11384);
not G12780 (W11383, I1329);
not G12781 (W11384, W13446);
not G12782 (W11385, W11387);
not G12783 (W11386, I1330);
not G12784 (W11387, W13447);
not G12785 (W11388, W11390);
not G12786 (W11389, I1331);
not G12787 (W11390, W13448);
not G12788 (W11391, W11393);
not G12789 (W11392, I1332);
not G12790 (W11393, W13449);
not G12791 (W11394, W11396);
not G12792 (W11395, I1333);
not G12793 (W11396, W13450);
not G12794 (W11397, W11399);
not G12795 (W11398, I1334);
not G12796 (W11399, W13451);
not G12797 (W11400, W11402);
not G12798 (W11401, I1335);
not G12799 (W11402, W13452);
not G12800 (W11403, W11405);
not G12801 (W11404, I1336);
not G12802 (W11405, W13453);
not G12803 (W11406, W11408);
not G12804 (W11407, I1337);
not G12805 (W11408, W13454);
not G12806 (W11409, W11411);
not G12807 (W11410, I1338);
not G12808 (W11411, W13455);
not G12809 (W11412, W11414);
not G12810 (W11413, I1339);
not G12811 (W11414, W13456);
not G12812 (W11415, W11417);
not G12813 (W11416, I1340);
not G12814 (W11417, W13457);
not G12815 (W11418, W11420);
not G12816 (W11419, I1341);
not G12817 (W11420, W13458);
not G12818 (W11421, W11423);
not G12819 (W11422, I1342);
not G12820 (W11423, W13459);
and G12821 (W11424, I1343, W13460);
and G12822 (W11425, W13461, W13462);
not G12823 (W11426, W13463);
not G12824 (W11427, W13464);
not G12825 (W11428, W13465);
and G12826 (W11429, W13466, W13467);
and G12827 (W11430, I1344, W13468);
and G12828 (W11431, I1345, W13469);
and G12829 (W11432, W13470, W13471);
and G12830 (W11433, W13472, W13473);
and G12831 (W11434, I1346, W13474);
and G12832 (W11435, I1347, W13475);
and G12833 (W11436, W13476, W13477);
and G12834 (W11437, W13478, W13479);
and G12835 (W11438, I1348, W13480);
and G12836 (W11439, I1349, W13481);
and G12837 (W11440, W13482, W13483);
and G12838 (W11441, W13484, W13485);
and G12839 (W11442, I1350, W13486);
and G12840 (W11443, I1351, W13487);
and G12841 (W11444, W13488, W13489);
and G12842 (W11445, W13490, W13491);
and G12843 (W11446, I1352, W13492);
and G12844 (W11447, W13493, W13494);
not G12845 (W11448, W11450);
not G12846 (W11449, I1353);
not G12847 (W11450, W13495);
not G12848 (W11451, W11453);
not G12849 (W11452, I1354);
not G12850 (W11453, W13496);
not G12851 (W11454, W11456);
not G12852 (W11455, I1355);
not G12853 (W11456, W13497);
not G12854 (W11457, W11459);
not G12855 (W11458, I1356);
not G12856 (W11459, W13498);
not G12857 (W11460, W11462);
not G12858 (W11461, I1357);
not G12859 (W11462, W13499);
not G12860 (W11463, W11465);
not G12861 (W11464, I1358);
not G12862 (W11465, W13500);
not G12863 (W11466, W11468);
not G12864 (W11467, I1359);
not G12865 (W11468, W13501);
not G12866 (W11469, W11471);
not G12867 (W11470, I1360);
not G12868 (W11471, W13502);
not G12869 (W11472, W11474);
not G12870 (W11473, I1361);
not G12871 (W11474, W13503);
nand G12872 (W11475, W11324, W11336, W13504);
not G12873 (W11476, W11478);
not G12874 (W11477, I1362);
not G12875 (W11478, W13505);
not G12876 (W11479, W11481);
not G12877 (W11480, I1363);
not G12878 (W11481, W13506);
not G12879 (W11482, W11484);
not G12880 (W11483, I1364);
not G12881 (W11484, W13507);
not G12882 (W11485, W13508);
not G12883 (W11486, W13509);
not G12884 (W11487, I209);
not G12885 (W11488, W11490);
nand G12886 (W11489, W13510, W13511);
not G12887 (W11490, W13512);
not G12888 (W11491, W11492);
not G12889 (W11492, W13513);
not G12890 (W11493, W11495);
nand G12891 (W11494, W13514, W13515);
not G12892 (W11495, W13516);
not G12893 (W11496, I200);
not G12894 (W11497, W11498);
not G12895 (W11498, W13517);
not G12896 (W11499, W13518);
not G12897 (W11500, W13519);
not G12898 (W11501, W13520);
not G12899 (W11502, W13521);
not G12900 (W11503, I223);
not G12901 (W11504, W11506);
not G12902 (W11505, I1365);
not G12903 (W11506, W13522);
not G12904 (W11507, I224);
not G12905 (W11508, W11510);
not G12906 (W11509, I1366);
not G12907 (W11510, W13523);
not G12908 (W11511, I225);
not G12909 (W11512, W11514);
not G12910 (W11513, I1367);
not G12911 (W11514, W13524);
not G12912 (W11515, I226);
not G12913 (W11516, W11518);
not G12914 (W11517, I1368);
not G12915 (W11518, W13525);
not G12916 (W11519, I227);
not G12917 (W11520, W11522);
not G12918 (W11521, I1369);
not G12919 (W11522, W13526);
not G12920 (W11523, I228);
not G12921 (W11524, W11526);
not G12922 (W11525, I1370);
not G12923 (W11526, W13527);
not G12924 (W11527, I229);
not G12925 (W11528, W11530);
not G12926 (W11529, I1371);
not G12927 (W11530, W13528);
not G12928 (W11531, I230);
not G12929 (W11532, W11534);
not G12930 (W11533, I1372);
not G12931 (W11534, W13529);
not G12932 (W11535, I201);
not G12933 (W11536, W11538);
not G12934 (W11537, I1373);
not G12935 (W11538, W13530);
not G12936 (W11539, I202);
not G12937 (W11540, W11542);
not G12938 (W11541, I1374);
not G12939 (W11542, W13531);
not G12940 (W11543, I203);
not G12941 (W11544, W11546);
not G12942 (W11545, I1375);
not G12943 (W11546, W13532);
not G12944 (W11547, I204);
not G12945 (W11548, W11550);
not G12946 (W11549, I1376);
not G12947 (W11550, W13533);
not G12948 (W11551, I205);
not G12949 (W11552, W11554);
not G12950 (W11553, I1377);
not G12951 (W11554, W13534);
not G12952 (W11555, I206);
not G12953 (W11556, W11558);
not G12954 (W11557, I1378);
not G12955 (W11558, W13535);
not G12956 (W11559, I207);
not G12957 (W11560, W11562);
not G12958 (W11561, I1379);
not G12959 (W11562, W13536);
not G12960 (W11563, I208);
not G12961 (W11564, W11566);
not G12962 (W11565, I1380);
not G12963 (W11566, W13537);
not G12964 (W11567, I210);
not G12965 (W11568, W11569);
not G12966 (W11569, W13538);
not G12967 (W11570, I211);
not G12968 (W11571, W11572);
not G12969 (W11572, W13539);
not G12970 (W11573, I212);
not G12971 (W11574, W11575);
not G12972 (W11575, W13540);
not G12973 (W11576, I213);
not G12974 (W11577, W11578);
not G12975 (W11578, W13541);
not G12976 (W11579, I214);
not G12977 (W11580, W11581);
not G12978 (W11581, W13542);
not G12979 (W11582, I215);
not G12980 (W11583, W11584);
not G12981 (W11584, W13543);
not G12982 (W11585, I216);
not G12983 (W11586, W11587);
not G12984 (W11587, W13544);
not G12985 (W11588, I217);
not G12986 (W11589, W11590);
not G12987 (W11590, W13545);
not G12988 (W11591, I247);
not G12989 (W11592, W11593);
not G12990 (W11593, W13546);
not G12991 (W11594, I248);
not G12992 (W11595, W11596);
not G12993 (W11596, W13547);
not G12994 (W11597, I249);
not G12995 (W11598, W11599);
not G12996 (W11599, W13548);
not G12997 (W11600, I250);
not G12998 (W11601, W11602);
not G12999 (W11602, W13549);
not G13000 (W11603, I251);
not G13001 (W11604, W11605);
not G13002 (W11605, W13550);
not G13003 (W11606, I252);
not G13004 (W11607, W11608);
not G13005 (W11608, W13551);
not G13006 (W11609, I253);
not G13007 (W11610, W11611);
not G13008 (W11611, W13552);
not G13009 (W11612, I254);
not G13010 (W11613, W11614);
not G13011 (W11614, W13553);
nand G13012 (W11615, I408, W11616);
nand G13013 (W11616, W13554, W13555);
nand G13014 (W11617, I409, W11618);
nand G13015 (W11618, W13556, W13557);
not G13016 (W11619, I218);
not G13017 (W11620, W13558);
and G13018 (W11621, W13559, W13560);
and G13019 (W11622, I1381, W13561);
and G13020 (W11623, W13562, W13563);
and G13021 (W11624, I1382, W13564);
and G13022 (W11625, I1383, W13565);
and G13023 (W11626, W13566, W13567);
and G13024 (W11627, I1384, W13568);
and G13025 (W11628, W13569, W13570);
and G13026 (W11629, W13566, I1381, W13571);
and G13027 (W11630, I1385, W13572);
and G13028 (W11631, W13573, W13574);
and G13029 (W11632, W13575, W13576);
and G13030 (W11633, I1386, W13577);
and G13031 (W11634, I1387, W13578);
and G13032 (W11635, W13579, W13580);
and G13033 (W11636, W13581, W13582);
and G13034 (W11637, I1388, W13583);
and G13035 (W11638, I1389, W13584);
and G13036 (W11639, W13585, W13586);
and G13037 (W11640, W13587, W13588);
and G13038 (W11641, I1390, W13589);
and G13039 (W11642, I1391, W13590);
and G13040 (W11643, W13591, W13592);
and G13041 (W11644, W13593, W13594);
not G13042 (W11645, W13595);
not G13043 (W11646, W13596);
not G13044 (W11647, W13597);
not G13045 (W11648, W13598);
not G13046 (W11649, I1392);
nand G13047 (W11650, W11649, W7919);
nand G13048 (W11651, W13599, W13600);
nand G13049 (W11652, W13601, W13600);
not G13050 (W11653, W13602);
not G13051 (W11654, I1393);
not G13052 (W11655, I1394);
nand G13053 (W11656, W11655, W7924);
nand G13054 (W11657, W13603, W13604);
nand G13055 (W11658, W13605, W13604);
not G13056 (W11659, W13606);
not G13057 (W11660, W13606);
not G13058 (W11661, W13606);
not G13059 (W11662, W13606);
not G13060 (W11663, W13606);
not G13061 (W11664, W13606);
not G13062 (W11665, W13606);
not G13063 (W11666, W13606);
not G13064 (W11667, W13606);
not G13065 (W11668, W13606);
not G13066 (W11669, W13606);
not G13067 (W11670, W13606);
not G13068 (W11671, W13606);
not G13069 (W11672, W13606);
not G13070 (W11673, W13606);
not G13071 (W11674, W13606);
not G13072 (W11675, W13606);
not G13073 (W11676, W13606);
not G13074 (W11677, W13607);
not G13075 (W11678, W11017);
not G13076 (W11679, W13607);
not G13077 (W11680, W10244);
not G13078 (W11681, W13607);
not G13079 (W11682, W9471);
not G13080 (W11683, W13607);
not G13081 (W11684, W8698);
nor G13082 (W11685, W13608, W13609);
not G13083 (W11686, W11015);
not G13084 (W11687, W11016);
not G13085 (W11688, W11017);
nor G13086 (W11689, W13610, W13611);
not G13087 (W11690, W11015);
not G13088 (W11691, W11016);
not G13089 (W11692, W11017);
nor G13090 (W11693, W13612, W13613);
not G13091 (W11694, W11015);
not G13092 (W11695, W11016);
not G13093 (W11696, W11017);
nor G13094 (W11697, W13612, W13614);
not G13095 (W11698, W11015);
not G13096 (W11699, W11016);
not G13097 (W11700, W11017);
nor G13098 (W11701, W13615, W13616);
not G13099 (W11702, W10242);
not G13100 (W11703, W10243);
not G13101 (W11704, W10244);
nor G13102 (W11705, W13617, W13618);
not G13103 (W11706, W10242);
not G13104 (W11707, W10243);
not G13105 (W11708, W10244);
nor G13106 (W11709, W13619, W13620);
not G13107 (W11710, W10242);
not G13108 (W11711, W10243);
not G13109 (W11712, W10244);
nor G13110 (W11713, W13619, W13621);
not G13111 (W11714, W10242);
not G13112 (W11715, W10243);
not G13113 (W11716, W10244);
nor G13114 (W11717, W13622, W13623);
not G13115 (W11718, W9469);
not G13116 (W11719, W9470);
not G13117 (W11720, W9471);
nor G13118 (W11721, W13624, W13625);
not G13119 (W11722, W9469);
not G13120 (W11723, W9470);
not G13121 (W11724, W9471);
nor G13122 (W11725, W13626, W13627);
not G13123 (W11726, W9469);
not G13124 (W11727, W9470);
not G13125 (W11728, W9471);
nor G13126 (W11729, W13626, W13628);
not G13127 (W11730, W9469);
not G13128 (W11731, W9470);
not G13129 (W11732, W9471);
nor G13130 (W11733, W13629, W13630);
not G13131 (W11734, W8696);
not G13132 (W11735, W8697);
not G13133 (W11736, W8698);
nor G13134 (W11737, W13631, W13632);
not G13135 (W11738, W8696);
not G13136 (W11739, W8697);
not G13137 (W11740, W8698);
nor G13138 (W11741, W13633, W13634);
not G13139 (W11742, W8696);
not G13140 (W11743, W8697);
not G13141 (W11744, W8698);
nor G13142 (W11745, W13633, W13635);
not G13143 (W11746, W8696);
not G13144 (W11747, W8697);
not G13145 (W11748, W8698);
not G13146 (W11749, I500);
not G13147 (W11750, W11751);
not G13148 (W11751, W13636);
not G13149 (W11752, I501);
not G13150 (W11753, W11754);
not G13151 (W11754, W13637);
not G13152 (W11755, W11757);
not G13153 (W11756, I502);
not G13154 (W11757, W13638);
not G13155 (W11758, W11760);
not G13156 (W11759, I503);
not G13157 (W11760, W13639);
and G13158 (W11761, W11874, I503, W11752);
not G13159 (W11762, W13640);
not G13160 (W11763, W13641);
not G13161 (W11764, W13642);
not G13162 (W11765, W13643);
nor G13163 (W11766, W13644, W13645, W13646);
nor G13164 (W11767, W13647, W13648);
not G13165 (W11768, W13649);
or G13166 (W11769, W5251, W13650);
or G13167 (W11770, W13651, W13652, W5253);
or G13168 (W11771, W13653, W13652, W13654);
not G13169 (W11772, W13655);
nor G13170 (W11773, W13656, W13657);
nor G13171 (W11774, W13658, W13659);
not G13172 (W11775, W13660);
or G13173 (W11776, W13661, W13653, W5253);
or G13174 (W11777, W13661, W13651, W13654);
not G13175 (W11778, W13662);
not G13176 (W11779, W13663);
not G13177 (W11780, W13664);
not G13178 (W11781, W13665);
not G13179 (W11782, W13666);
not G13180 (W11783, W13667);
not G13181 (W11784, W13668);
not G13182 (W11785, W13669);
not G13183 (W11786, W13670);
not G13184 (W11787, W13671);
not G13185 (W11788, W11018);
not G13186 (W11789, W8243);
not G13187 (W11790, W13672);
nor G13188 (W11791, W13673, W13674, W13675);
nor G13189 (W11792, W13676, W13677, W13678);
nor G13190 (W11793, W13679, W13680, W13681);
nor G13191 (W11794, W13682, W13683);
not G13192 (W11795, W13684);
or G13193 (W11796, W4976, W13685);
or G13194 (W11797, W13686, W13687, W4978);
or G13195 (W11798, W13688, W13687, W13689);
not G13196 (W11799, W13690);
nor G13197 (W11800, W13691, W13692);
nor G13198 (W11801, W13693, W13694);
not G13199 (W11802, W13695);
or G13200 (W11803, W13696, W13688, W4978);
or G13201 (W11804, W13696, W13686, W13689);
not G13202 (W11805, W13697);
not G13203 (W11806, W13698);
not G13204 (W11807, W13699);
not G13205 (W11808, W13700);
not G13206 (W11809, W13701);
not G13207 (W11810, W13702);
not G13208 (W11811, W13703);
not G13209 (W11812, W13704);
not G13210 (W11813, W13705);
not G13211 (W11814, W13706);
not G13212 (W11815, W10245);
not G13213 (W11816, W8286);
nor G13214 (W11817, W13707, W13708, W13709);
nor G13215 (W11818, W13710, W13711, W13712);
nor G13216 (W11819, W13713, W13714, W13715);
nor G13217 (W11820, W13716, W13717);
not G13218 (W11821, W13718);
or G13219 (W11822, W4701, W13719);
or G13220 (W11823, W13720, W13721, W4703);
or G13221 (W11824, W13722, W13721, W13723);
not G13222 (W11825, W13724);
nor G13223 (W11826, W13725, W13726);
nor G13224 (W11827, W13727, W13728);
not G13225 (W11828, W13729);
or G13226 (W11829, W13730, W13722, W4703);
or G13227 (W11830, W13730, W13720, W13723);
not G13228 (W11831, W13731);
not G13229 (W11832, W13732);
not G13230 (W11833, W13733);
not G13231 (W11834, W13734);
not G13232 (W11835, W13735);
not G13233 (W11836, W13736);
not G13234 (W11837, W13737);
not G13235 (W11838, W13738);
not G13236 (W11839, W13739);
not G13237 (W11840, W13740);
not G13238 (W11841, W9472);
not G13239 (W11842, W8329);
nor G13240 (W11843, W13741, W13742, W13743);
nor G13241 (W11844, W13744, W13745, W13746);
nor G13242 (W11845, W13747, W13748, W13749);
nor G13243 (W11846, W13750, W13751);
not G13244 (W11847, W13752);
or G13245 (W11848, W4426, W13753);
or G13246 (W11849, W13754, W13755, W4428);
or G13247 (W11850, W13756, W13755, W13757);
not G13248 (W11851, W13758);
nor G13249 (W11852, W13759, W13760);
nor G13250 (W11853, W13761, W13762);
not G13251 (W11854, W13763);
or G13252 (W11855, W13764, W13756, W4428);
or G13253 (W11856, W13764, W13754, W13757);
not G13254 (W11857, W13765);
not G13255 (W11858, W13766);
not G13256 (W11859, W13767);
not G13257 (W11860, W13768);
not G13258 (W11861, W13769);
not G13259 (W11862, W13770);
not G13260 (W11863, W13771);
not G13261 (W11864, W13772);
not G13262 (W11865, W13773);
not G13263 (W11866, W13774);
not G13264 (W11867, W8699);
not G13265 (W11868, W8372);
nor G13266 (W11869, W13775, W13776, W13777);
nor G13267 (W11870, W13778, W13779, W13780);
not G13268 (W11871, W11873);
not G13269 (W11872, I556);
not G13270 (W11873, W13781);
and G13271 (W11874, W13782, W13783);
and G13272 (W11875, I1395, W13784);
and G13273 (W11876, W13785, W13786);
not G13274 (W11877, W8376);
and G13275 (W11878, W13787, W13788);
and G13276 (W11879, I1396, W13789);
not G13277 (W11880, W5837);
not G13278 (W11881, W11883);
not G13279 (W11882, I557);
not G13280 (W11883, W13790);
not G13281 (W11884, I558);
not G13282 (W11885, W11886);
not G13283 (W11886, W13791);
not G13284 (W11887, W11889);
not G13285 (W11888, I559);
not G13286 (W11889, W13792);
not G13287 (W11890, I560);
not G13288 (W11891, W11892);
not G13289 (W11892, W13793);
not G13290 (W11893, I257);
not G13291 (W11894, W13794);
nor G13292 (W11895, W13795, W13796);
not G13293 (W11896, W11898);
nor G13294 (W11897, W13797, W13798);
not G13295 (W11898, W13799);
nor G13296 (W11899, W13795, W13796);
not G13297 (W11900, W11902);
nor G13298 (W11901, W13800, W13801);
not G13299 (W11902, W13802);
nor G13300 (W11903, W13803, W13796);
not G13301 (W11904, W11906);
nor G13302 (W11905, W13804, W13805);
not G13303 (W11906, W13806);
nor G13304 (W11907, W13803, W13796);
not G13305 (W11908, W11910);
nor G13306 (W11909, W13807, W13808);
not G13307 (W11910, W13809);
nor G13308 (W11911, W13810, W13796);
not G13309 (W11912, W11914);
nor G13310 (W11913, W13811, W13812);
not G13311 (W11914, W13813);
nor G13312 (W11915, W11867, W11917);
and G13313 (W11916, W13814, W13815, W13816);
not G13314 (W11917, W8701);
nand G13315 (W11918, W13817, W13818);
nand G13316 (W11919, W13819, W13820);
nor G13317 (W11920, W13821, W13796);
not G13318 (W11921, W11923);
nor G13319 (W11922, W13822, W13823);
not G13320 (W11923, W13824);
nor G13321 (W11924, W13825, W13796);
not G13322 (W11925, W11927);
nor G13323 (W11926, W13826, W13827);
not G13324 (W11927, W13828);
nor G13325 (W11928, W13825, W13796);
not G13326 (W11929, W11931);
nor G13327 (W11930, W13829, W13830);
not G13328 (W11931, W13831);
not G13329 (W11932, I603);
not G13330 (W11933, W13832);
not G13331 (W11934, W13833);
not G13332 (W11935, W13834);
nor G13333 (W11936, W13835, W13836, W13837);
not G13334 (W11937, W13838);
not G13335 (W11938, W13839);
not G13336 (W11939, W13840);
not G13337 (W11940, W8373);
not G13338 (W11941, W13841);
not G13339 (W11942, W13842);
not G13340 (W11943, W13843);
not G13341 (W11944, W11866);
not G13342 (W11945, W13844);
not G13343 (W11946, W13845);
not G13344 (W11947, W13846);
not G13345 (W11948, W13847);
not G13346 (W11949, W13848);
not G13347 (W11950, W13849);
not G13348 (W11951, W13850);
not G13349 (W11952, W13851);
not G13350 (W11953, W13852);
not G13351 (W11954, W13853);
not G13352 (W11955, W13854);
not G13353 (W11956, W13855);
not G13354 (W11957, W13856);
not G13355 (W11958, W13857);
not G13356 (W11959, W13858);
not G13357 (W11960, W13859);
not G13358 (W11961, W13860);
not G13359 (W11962, W13861);
not G13360 (W11963, W13862);
not G13361 (W11964, W13863);
not G13362 (W11965, W13864);
not G13363 (W11966, W13865);
not G13364 (W11967, W13866);
not G13365 (W11968, W13867);
not G13366 (W11969, W13868);
not G13367 (W11970, W13869);
not G13368 (W11971, W13870);
not G13369 (W11972, W13871);
not G13370 (W11973, W13872);
not G13371 (W11974, W13873);
not G13372 (W11975, W13874);
not G13373 (W11976, W13875);
not G13374 (W11977, W13876);
not G13375 (W11978, W11980);
not G13376 (W11979, I260);
not G13377 (W11980, W13877);
not G13378 (W11981, I2);
not G13379 (W11982, I261);
not G13380 (W11983, W11984);
not G13381 (W11984, W13878);
not G13382 (W11985, W11987);
not G13383 (W11986, I262);
not G13384 (W11987, W13879);
not G13385 (W11988, I263);
not G13386 (W11989, W11990);
not G13387 (W11990, W13880);
not G13388 (W11991, W11993);
not G13389 (W11992, I264);
not G13390 (W11993, W13881);
not G13391 (W11994, I265);
not G13392 (W11995, W11996);
not G13393 (W11996, W13882);
not G13394 (W11997, W11999);
not G13395 (W11998, I266);
not G13396 (W11999, W13883);
not G13397 (W12000, I267);
not G13398 (W12001, W12002);
not G13399 (W12002, W13884);
not G13400 (W12003, W12005);
not G13401 (W12004, I268);
not G13402 (W12005, W13885);
not G13403 (W12006, I269);
not G13404 (W12007, W12008);
not G13405 (W12008, W13886);
not G13406 (W12009, W13643);
and G13407 (W12010, I4, W13887);
and G13408 (W12011, W13888, W13889);
not G13409 (W12012, W13890);
and G13410 (W12013, I1397, W13891);
and G13411 (W12014, W13892, W13893);
not G13412 (W12015, W13890);
and G13413 (W12016, I1398, W13894);
and G13414 (W12017, W13895, W13896);
not G13415 (W12018, W13890);
and G13416 (W12019, I1399, W13897);
and G13417 (W12020, W13898, W13899);
not G13418 (W12021, W13890);
and G13419 (W12022, I1400, W13900);
and G13420 (W12023, W13901, W13902);
not G13421 (W12024, W13890);
not G13422 (W12025, W13903);
not G13423 (W12026, W8698);
not G13424 (W12027, W8696);
not G13425 (W12028, W8697);
not G13426 (W12029, W13904);
not G13427 (W12030, W13905);
not G13428 (W12031, W13906);
not G13429 (W12032, W13907);
not G13430 (W12033, W13908);
not G13431 (W12034, W13905);
not G13432 (W12035, W13906);
not G13433 (W12036, W13907);
and G13434 (W12037, I1401, W13909);
and G13435 (W12038, W12446, W13910);
not G13436 (W12039, I219);
not G13437 (W12040, W13911);
not G13438 (W12041, W13905);
not G13439 (W12042, W13906);
not G13440 (W12043, W13907);
not G13441 (W12044, W13912);
not G13442 (W12045, W13913);
not G13443 (W12046, W13914);
not G13444 (W12047, W13915);
and G13445 (W12048, W8697, W8661);
and G13446 (W12049, W8698, W8658);
and G13447 (W12050, W8696, W8654);
not G13448 (W12051, W4560);
not G13449 (W12052, W13913);
not G13450 (W12053, W13914);
not G13451 (W12054, W13915);
and G13452 (W12055, W8697, W8672);
and G13453 (W12056, W8698, W8669);
and G13454 (W12057, W8696, W8665);
not G13455 (W12058, W13916);
not G13456 (W12059, W13913);
not G13457 (W12060, W13914);
not G13458 (W12061, W13915);
not G13459 (W12062, W13917);
not G13460 (W12063, W13913);
not G13461 (W12064, W13914);
not G13462 (W12065, W13915);
and G13463 (W12066, W8697, W8693);
and G13464 (W12067, W8698, W8690);
and G13465 (W12068, W8696, W8686);
not G13466 (W12069, W13918);
not G13467 (W12070, W13913);
not G13468 (W12071, W13914);
not G13469 (W12072, W13915);
not G13470 (W12073, I21);
not G13471 (W12074, I20);
not G13472 (W12075, I1402);
not G13473 (W12076, W8698);
not G13474 (W12077, W8698);
and G13475 (W12078, W13919, W13920);
and G13476 (W12079, W13921, W13922);
not G13477 (W12080, W13923);
and G13478 (W12081, W13924, W13925);
and G13479 (W12082, W13926, W13927);
not G13480 (W12083, W13923);
and G13481 (W12084, I1403, W13928);
and G13482 (W12085, W13929, W13930);
not G13483 (W12086, W13923);
and G13484 (W12087, I1404, W13931);
and G13485 (W12088, W13932, W13933);
not G13486 (W12089, W13923);
and G13487 (W12090, I1405, W13934);
and G13488 (W12091, W13935, W13936);
not G13489 (W12092, W13923);
and G13490 (W12093, I1406, W13937);
and G13491 (W12094, W13938, W13939);
not G13492 (W12095, W13923);
and G13493 (W12096, I638, W13940);
and G13494 (W12097, W13941, W13942);
not G13495 (W12098, W13943);
not G13496 (W12099, W13944);
not G13497 (W12100, W13945);
not G13498 (W12101, W13946);
not G13499 (W12102, W13947);
nor G13500 (W12103, W13948, W13949);
not G13501 (W12104, W13950);
not G13502 (W12105, W13951);
not G13503 (W12106, W9107);
nor G13504 (W12107, W13952, W13953);
not G13505 (W12108, W13950);
not G13506 (W12109, W13951);
not G13507 (W12110, W9107);
nor G13508 (W12111, W13954, W13955);
not G13509 (W12112, W13950);
not G13510 (W12113, W13951);
not G13511 (W12114, W9107);
nor G13512 (W12115, W13956, W13957);
not G13513 (W12116, W13950);
not G13514 (W12117, W13951);
not G13515 (W12118, W9107);
nor G13516 (W12119, W13958, W13959);
not G13517 (W12120, W9107);
not G13518 (W12121, W13950);
not G13519 (W12122, W13951);
nor G13520 (W12123, W13960, W13961);
not G13521 (W12124, W13951);
not G13522 (W12125, W9107);
not G13523 (W12126, W13950);
nor G13524 (W12127, W13962, W13963);
not G13525 (W12128, W13950);
not G13526 (W12129, W13951);
not G13527 (W12130, W9107);
nor G13528 (W12131, W13964, W13965);
not G13529 (W12132, W13950);
not G13530 (W12133, W13951);
not G13531 (W12134, W9107);
nor G13532 (W12135, W13966, W13967);
not G13533 (W12136, W13950);
not G13534 (W12137, W13951);
not G13535 (W12138, W9107);
nor G13536 (W12139, W13968, W13969);
not G13537 (W12140, W13950);
not G13538 (W12141, W13951);
not G13539 (W12142, W9107);
nor G13540 (W12143, W13970, W13971);
not G13541 (W12144, W12210);
not G13542 (W12145, W12211);
not G13543 (W12146, W12212);
nor G13544 (W12147, W13970, W13972);
not G13545 (W12148, W12210);
not G13546 (W12149, W12211);
not G13547 (W12150, W12212);
nor G13548 (W12151, W13970, W13973);
not G13549 (W12152, W12210);
not G13550 (W12153, W12211);
not G13551 (W12154, W12212);
nor G13552 (W12155, W13974, W13975);
not G13553 (W12156, W13976);
not G13554 (W12157, W13977);
not G13555 (W12158, W13978);
not G13556 (W12159, W13979);
nand G13557 (W12160, W13980, W13981);
nor G13558 (W12161, W13982, W13983, W13984);
and G13559 (W12162, W13985, W13986);
nor G13560 (W12163, W13987, W13988, W13989);
nor G13561 (W12164, W13990, W13991);
not G13562 (W12165, W13992);
or G13563 (W12166, W4565, W13993);
or G13564 (W12167, W13994, W13995, W4573);
or G13565 (W12168, W13996, W13995, W13997);
not G13566 (W12169, W13998);
nor G13567 (W12170, W13999, W14000);
nor G13568 (W12171, W14001, W14002);
not G13569 (W12172, W14003);
or G13570 (W12173, W14004, W13996, W4573);
or G13571 (W12174, W14004, W13994, W13997);
not G13572 (W12175, W14005);
not G13573 (W12176, W14006);
not G13574 (W12177, W14007);
not G13575 (W12178, W14008);
not G13576 (W12179, W14009);
not G13577 (W12180, W14010);
not G13578 (W12181, W14011);
not G13579 (W12182, W14012);
not G13580 (W12183, W14013);
nand G13581 (W12184, W14014, W14015);
not G13582 (W12185, W12210);
not G13583 (W12186, W12211);
not G13584 (W12187, W12212);
not G13585 (W12188, I1407);
not G13586 (W12189, W14016);
nor G13587 (W12190, W14017, W14018);
not G13588 (W12191, W14019);
not G13589 (W12192, W14020);
not G13590 (W12193, W14021);
not G13591 (W12194, W14022);
not G13592 (W12195, W12212);
not G13593 (W12196, W12210);
not G13594 (W12197, W12211);
nand G13595 (W12198, W14023, W14024);
not G13596 (W12199, W12210);
not G13597 (W12200, W12211);
not G13598 (W12201, W12212);
nand G13599 (W12202, W14025, W14026);
not G13600 (W12203, W12210);
not G13601 (W12204, W12211);
not G13602 (W12205, W12212);
not G13603 (W12206, W14027);
not G13604 (W12207, W14028);
not G13605 (W12208, W14029);
not G13606 (W12209, W14030);
not G13607 (W12210, W14031);
not G13608 (W12211, W14032);
not G13609 (W12212, W14033);
not G13610 (W12213, I225);
not G13611 (W12214, W14034);
not G13612 (W12215, I226);
not G13613 (W12216, W14035);
not G13614 (W12217, I227);
not G13615 (W12218, W14036);
not G13616 (W12219, I228);
not G13617 (W12220, W14037);
not G13618 (W12221, I229);
not G13619 (W12222, W14038);
not G13620 (W12223, I230);
not G13621 (W12224, W14039);
nor G13622 (W12225, W14040, W14041, W14042);
not G13623 (W12226, W14043);
not G13624 (W12227, I223);
not G13625 (W12228, W14044);
nor G13626 (W12229, W14045, W14046, W14047);
not G13627 (W12230, W14048);
not G13628 (W12231, I224);
not G13629 (W12232, W14049);
not G13630 (W12233, W14050);
not G13631 (W12234, W14051);
not G13632 (W12235, W14052);
not G13633 (W12236, W14053);
not G13634 (W12237, W14054);
not G13635 (W12238, W14055);
not G13636 (W12239, W14056);
not G13637 (W12240, W14057);
not G13638 (W12241, W14058);
not G13639 (W12242, W14059);
not G13640 (W12243, W14060);
not G13641 (W12244, W14061);
not G13642 (W12245, W14062);
not G13643 (W12246, W14063);
not G13644 (W12247, W14064);
not G13645 (W12248, W14065);
not G13646 (W12249, W14066);
not G13647 (W12250, W14067);
not G13648 (W12251, W14068);
not G13649 (W12252, W14069);
not G13650 (W12253, W12255);
not G13651 (W12254, I740);
not G13652 (W12255, W14070);
not G13653 (W12256, I1408);
not G13654 (W12257, I1409);
not G13655 (W12258, W13986);
not G13656 (W12259, I741);
not G13657 (W12260, W12261);
not G13658 (W12261, W14071);
not G13659 (W12262, W12264);
not G13660 (W12263, I742);
not G13661 (W12264, W14072);
not G13662 (W12265, I743);
not G13663 (W12266, W12267);
not G13664 (W12267, W14073);
not G13665 (W12268, W12270);
not G13666 (W12269, I744);
not G13667 (W12270, W14074);
not G13668 (W12271, I745);
not G13669 (W12272, W12273);
not G13670 (W12273, W14075);
not G13671 (W12274, W12276);
not G13672 (W12275, I746);
not G13673 (W12276, W14076);
not G13674 (W12277, I747);
not G13675 (W12278, W12279);
not G13676 (W12279, W14077);
not G13677 (W12280, W12282);
not G13678 (W12281, I748);
not G13679 (W12282, W14078);
not G13680 (W12283, I749);
not G13681 (W12284, W12285);
not G13682 (W12285, W14079);
and G13683 (W12286, W9033, W9041, W9005, W9009);
and G13684 (W12287, W9013, W9017, W9021, W9025);
not G13685 (W12288, W14080);
not G13686 (W12289, W14081);
not G13687 (W12290, W14082);
not G13688 (W12291, W14083);
not G13689 (W12292, W14084);
not G13690 (W12293, W14085);
not G13691 (W12294, W14086);
not G13692 (W12295, W14087);
not G13693 (W12296, W14088);
nor G13694 (W12297, W9017, W9021);
not G13695 (W12298, W14089);
not G13696 (W12299, W14090);
not G13697 (W12300, W14091);
nor G13698 (W12301, W14092, W14093);
not G13699 (W12302, W12304);
nor G13700 (W12303, W14094, W14095);
not G13701 (W12304, W14096);
nor G13702 (W12305, W14092, W14093);
not G13703 (W12306, W12308);
nor G13704 (W12307, W14097, W14098);
not G13705 (W12308, W14099);
nor G13706 (W12309, W14100, W14093);
not G13707 (W12310, W12312);
nor G13708 (W12311, W14101, W14102);
not G13709 (W12312, W14103);
nor G13710 (W12313, W14100, W14093);
not G13711 (W12314, W12316);
nor G13712 (W12315, W14104, W14105);
not G13713 (W12316, W14106);
nor G13714 (W12317, W14107, W14093);
not G13715 (W12318, W12320);
nor G13716 (W12319, W14108, W14109);
not G13717 (W12320, W14110);
nor G13718 (W12321, W11841, W12323);
and G13719 (W12322, W14111, W14112, W14113);
not G13720 (W12323, W9474);
nand G13721 (W12324, W14114, W14115);
nand G13722 (W12325, W14116, W14117);
nor G13723 (W12326, W14118, W14093);
not G13724 (W12327, W12329);
nor G13725 (W12328, W14119, W14120);
not G13726 (W12329, W14121);
nor G13727 (W12330, W14122, W14093);
not G13728 (W12331, W12333);
nor G13729 (W12332, W14123, W14124);
not G13730 (W12333, W14125);
nor G13731 (W12334, W14122, W14093);
not G13732 (W12335, W12337);
nor G13733 (W12336, W14126, W14127);
not G13734 (W12337, W14128);
not G13735 (W12338, I804);
not G13736 (W12339, W14129);
not G13737 (W12340, W14130);
not G13738 (W12341, W14131);
nor G13739 (W12342, W14132, W14133, W14134);
not G13740 (W12343, W14135);
not G13741 (W12344, W14136);
not G13742 (W12345, W14137);
not G13743 (W12346, W8330);
not G13744 (W12347, W14138);
not G13745 (W12348, W14139);
not G13746 (W12349, W14140);
not G13747 (W12350, W11840);
not G13748 (W12351, W14141);
not G13749 (W12352, W14142);
not G13750 (W12353, W14143);
not G13751 (W12354, W14144);
not G13752 (W12355, W14145);
not G13753 (W12356, W14146);
not G13754 (W12357, W14147);
not G13755 (W12358, W14148);
not G13756 (W12359, W14149);
not G13757 (W12360, W14150);
not G13758 (W12361, W14151);
not G13759 (W12362, W14152);
not G13760 (W12363, W14153);
not G13761 (W12364, W14154);
not G13762 (W12365, W14155);
not G13763 (W12366, W14156);
not G13764 (W12367, W14157);
not G13765 (W12368, W14158);
not G13766 (W12369, W14159);
not G13767 (W12370, W14160);
not G13768 (W12371, W14161);
not G13769 (W12372, W14162);
not G13770 (W12373, W14163);
not G13771 (W12374, W14164);
not G13772 (W12375, W14165);
not G13773 (W12376, W14166);
not G13774 (W12377, W14167);
not G13775 (W12378, W14168);
not G13776 (W12379, W14169);
not G13777 (W12380, W14170);
not G13778 (W12381, W14171);
not G13779 (W12382, W14172);
not G13780 (W12383, W14173);
not G13781 (W12384, W12386);
not G13782 (W12385, I296);
not G13783 (W12386, W14174);
not G13784 (W12387, I51);
not G13785 (W12388, I297);
not G13786 (W12389, W12390);
not G13787 (W12390, W14175);
not G13788 (W12391, W12393);
not G13789 (W12392, I298);
not G13790 (W12393, W14176);
not G13791 (W12394, I299);
not G13792 (W12395, W12396);
not G13793 (W12396, W14177);
not G13794 (W12397, W12399);
not G13795 (W12398, I300);
not G13796 (W12399, W14178);
not G13797 (W12400, I301);
not G13798 (W12401, W12402);
not G13799 (W12402, W14179);
not G13800 (W12403, W12405);
not G13801 (W12404, I302);
not G13802 (W12405, W14180);
not G13803 (W12406, I303);
not G13804 (W12407, W12408);
not G13805 (W12408, W14181);
not G13806 (W12409, W12411);
not G13807 (W12410, I304);
not G13808 (W12411, W14182);
not G13809 (W12412, I305);
not G13810 (W12413, W12414);
not G13811 (W12414, W14183);
not G13812 (W12415, W13642);
and G13813 (W12416, I53, W14184);
and G13814 (W12417, W14185, W14186);
not G13815 (W12418, W14187);
and G13816 (W12419, I1410, W14188);
and G13817 (W12420, W14189, W14190);
not G13818 (W12421, W14187);
and G13819 (W12422, I1411, W14191);
and G13820 (W12423, W14192, W14193);
not G13821 (W12424, W14187);
and G13822 (W12425, I1412, W14194);
and G13823 (W12426, W14195, W14196);
not G13824 (W12427, W14187);
and G13825 (W12428, I1413, W14197);
and G13826 (W12429, W14198, W14199);
not G13827 (W12430, W14187);
not G13828 (W12431, W14200);
not G13829 (W12432, W9471);
not G13830 (W12433, W9469);
not G13831 (W12434, W9470);
not G13832 (W12435, W14201);
not G13833 (W12436, W13905);
not G13834 (W12437, W13906);
not G13835 (W12438, W13907);
not G13836 (W12439, W14202);
not G13837 (W12440, W13905);
not G13838 (W12441, W13906);
not G13839 (W12442, W13907);
and G13840 (W12443, I1414, W14203);
and G13841 (W12444, W12852, W14204);
not G13842 (W12445, I220);
not G13843 (W12446, W14205);
not G13844 (W12447, W13905);
not G13845 (W12448, W13906);
not G13846 (W12449, W13907);
not G13847 (W12450, W14206);
not G13848 (W12451, W14207);
not G13849 (W12452, W14208);
not G13850 (W12453, W14209);
and G13851 (W12454, W9470, W9434);
and G13852 (W12455, W9471, W9431);
and G13853 (W12456, W9469, W9427);
not G13854 (W12457, W4835);
not G13855 (W12458, W14207);
not G13856 (W12459, W14208);
not G13857 (W12460, W14209);
and G13858 (W12461, W9470, W9445);
and G13859 (W12462, W9471, W9442);
and G13860 (W12463, W9469, W9438);
not G13861 (W12464, W14210);
not G13862 (W12465, W14207);
not G13863 (W12466, W14208);
not G13864 (W12467, W14209);
not G13865 (W12468, W14211);
not G13866 (W12469, W14207);
not G13867 (W12470, W14208);
not G13868 (W12471, W14209);
and G13869 (W12472, W9470, W9466);
and G13870 (W12473, W9471, W9463);
and G13871 (W12474, W9469, W9459);
not G13872 (W12475, W14212);
not G13873 (W12476, W14207);
not G13874 (W12477, W14208);
not G13875 (W12478, W14209);
not G13876 (W12479, I70);
not G13877 (W12480, I69);
not G13878 (W12481, I1415);
not G13879 (W12482, W9471);
not G13880 (W12483, W9471);
and G13881 (W12484, W14213, W14214);
and G13882 (W12485, W14215, W14216);
not G13883 (W12486, W14217);
and G13884 (W12487, W14218, W14219);
and G13885 (W12488, W14220, W14221);
not G13886 (W12489, W14217);
and G13887 (W12490, I1416, W14222);
and G13888 (W12491, W14223, W14224);
not G13889 (W12492, W14217);
and G13890 (W12493, I1417, W14225);
and G13891 (W12494, W14226, W14227);
not G13892 (W12495, W14217);
and G13893 (W12496, I1418, W14228);
and G13894 (W12497, W14229, W14230);
not G13895 (W12498, W14217);
and G13896 (W12499, I1419, W14231);
and G13897 (W12500, W14232, W14233);
not G13898 (W12501, W14217);
and G13899 (W12502, I839, W14234);
and G13900 (W12503, W14235, W14236);
not G13901 (W12504, W14237);
not G13902 (W12505, W14238);
not G13903 (W12506, W14239);
not G13904 (W12507, W14240);
not G13905 (W12508, W14241);
nor G13906 (W12509, W14242, W14243);
not G13907 (W12510, W14244);
not G13908 (W12511, W14245);
not G13909 (W12512, W9880);
nor G13910 (W12513, W14246, W14247);
not G13911 (W12514, W14244);
not G13912 (W12515, W14245);
not G13913 (W12516, W9880);
nor G13914 (W12517, W14248, W14249);
not G13915 (W12518, W14244);
not G13916 (W12519, W14245);
not G13917 (W12520, W9880);
nor G13918 (W12521, W14250, W14251);
not G13919 (W12522, W14244);
not G13920 (W12523, W14245);
not G13921 (W12524, W9880);
nor G13922 (W12525, W14252, W14253);
not G13923 (W12526, W14244);
not G13924 (W12527, W14245);
not G13925 (W12528, W9880);
nor G13926 (W12529, W14254, W14255);
not G13927 (W12530, W9880);
not G13928 (W12531, W14244);
not G13929 (W12532, W14245);
nor G13930 (W12533, W14256, W14257);
not G13931 (W12534, W14245);
not G13932 (W12535, W9880);
not G13933 (W12536, W14244);
nor G13934 (W12537, W14258, W14259);
not G13935 (W12538, W14245);
not G13936 (W12539, W9880);
not G13937 (W12540, W14244);
nor G13938 (W12541, W14260, W14261);
not G13939 (W12542, W14244);
not G13940 (W12543, W14245);
not G13941 (W12544, W9880);
nor G13942 (W12545, W14262, W14263);
not G13943 (W12546, W14244);
not G13944 (W12547, W14245);
not G13945 (W12548, W9880);
nor G13946 (W12549, W14264, W14265);
not G13947 (W12550, W12616);
not G13948 (W12551, W12617);
not G13949 (W12552, W12618);
nor G13950 (W12553, W14264, W14266);
not G13951 (W12554, W12616);
not G13952 (W12555, W12617);
not G13953 (W12556, W12618);
nor G13954 (W12557, W14264, W14267);
not G13955 (W12558, W12616);
not G13956 (W12559, W12617);
not G13957 (W12560, W12618);
nor G13958 (W12561, W14268, W14269);
not G13959 (W12562, W14270);
not G13960 (W12563, W14271);
not G13961 (W12564, W14272);
not G13962 (W12565, W14273);
nand G13963 (W12566, W14274, W14275);
nor G13964 (W12567, W14276, W14277, W14278);
and G13965 (W12568, W14279, W13986);
nor G13966 (W12569, W14280, W14281, W14282);
nor G13967 (W12570, W14283, W14284);
not G13968 (W12571, W14285);
or G13969 (W12572, W4840, W14286);
or G13970 (W12573, W14287, W14288, W4848);
or G13971 (W12574, W14289, W14288, W14290);
not G13972 (W12575, W14291);
nor G13973 (W12576, W14292, W14293);
nor G13974 (W12577, W14294, W14295);
not G13975 (W12578, W14296);
or G13976 (W12579, W14297, W14289, W4848);
or G13977 (W12580, W14297, W14287, W14290);
not G13978 (W12581, W14298);
not G13979 (W12582, W14299);
not G13980 (W12583, W14300);
not G13981 (W12584, W14301);
not G13982 (W12585, W14302);
not G13983 (W12586, W14303);
not G13984 (W12587, W14304);
not G13985 (W12588, W14305);
not G13986 (W12589, W14306);
nand G13987 (W12590, W14307, W14308);
not G13988 (W12591, W12616);
not G13989 (W12592, W12617);
not G13990 (W12593, W12618);
not G13991 (W12594, I1420);
not G13992 (W12595, W14309);
nor G13993 (W12596, W14310, W14311);
not G13994 (W12597, W14312);
not G13995 (W12598, W14313);
not G13996 (W12599, W14314);
not G13997 (W12600, W14315);
not G13998 (W12601, W12618);
not G13999 (W12602, W12616);
not G14000 (W12603, W12617);
nand G14001 (W12604, W14316, W14317);
not G14002 (W12605, W12616);
not G14003 (W12606, W12617);
not G14004 (W12607, W12618);
nand G14005 (W12608, W14318, W14319);
not G14006 (W12609, W12616);
not G14007 (W12610, W12617);
not G14008 (W12611, W12618);
not G14009 (W12612, W14320);
not G14010 (W12613, W14321);
not G14011 (W12614, W14322);
not G14012 (W12615, W14323);
not G14013 (W12616, W14324);
not G14014 (W12617, W14325);
not G14015 (W12618, W14326);
not G14016 (W12619, I249);
not G14017 (W12620, W14327);
not G14018 (W12621, I250);
not G14019 (W12622, W14328);
not G14020 (W12623, I251);
not G14021 (W12624, W14329);
not G14022 (W12625, I252);
not G14023 (W12626, W14330);
not G14024 (W12627, I253);
not G14025 (W12628, W14331);
not G14026 (W12629, I254);
not G14027 (W12630, W14332);
nor G14028 (W12631, W14333, W14334, W14335);
not G14029 (W12632, W14336);
not G14030 (W12633, I247);
not G14031 (W12634, W14337);
nor G14032 (W12635, W14338, W14339, W14340);
not G14033 (W12636, W14341);
not G14034 (W12637, I248);
not G14035 (W12638, W14342);
not G14036 (W12639, W14343);
not G14037 (W12640, W14344);
not G14038 (W12641, W14345);
not G14039 (W12642, W14346);
not G14040 (W12643, W14347);
not G14041 (W12644, W14348);
not G14042 (W12645, W14349);
not G14043 (W12646, W14350);
not G14044 (W12647, W14351);
not G14045 (W12648, W14352);
not G14046 (W12649, W14353);
not G14047 (W12650, W14354);
not G14048 (W12651, W14355);
not G14049 (W12652, W14356);
not G14050 (W12653, W14357);
not G14051 (W12654, W14358);
not G14052 (W12655, W14359);
not G14053 (W12656, W14360);
not G14054 (W12657, W14361);
not G14055 (W12658, W14362);
not G14056 (W12659, W12661);
not G14057 (W12660, I941);
not G14058 (W12661, W14363);
not G14059 (W12662, I1421);
not G14060 (W12663, I1422);
not G14061 (W12664, W13986);
not G14062 (W12665, I942);
not G14063 (W12666, W12667);
not G14064 (W12667, W14364);
not G14065 (W12668, W12670);
not G14066 (W12669, I943);
not G14067 (W12670, W14365);
not G14068 (W12671, I944);
not G14069 (W12672, W12673);
not G14070 (W12673, W14366);
not G14071 (W12674, W12676);
not G14072 (W12675, I945);
not G14073 (W12676, W14367);
not G14074 (W12677, I946);
not G14075 (W12678, W12679);
not G14076 (W12679, W14368);
not G14077 (W12680, W12682);
not G14078 (W12681, I947);
not G14079 (W12682, W14369);
not G14080 (W12683, I948);
not G14081 (W12684, W12685);
not G14082 (W12685, W14370);
not G14083 (W12686, W12688);
not G14084 (W12687, I949);
not G14085 (W12688, W14371);
not G14086 (W12689, I950);
not G14087 (W12690, W12691);
not G14088 (W12691, W14372);
and G14089 (W12692, W9806, W9814, W9778, W9782);
and G14090 (W12693, W9786, W9790, W9794, W9798);
not G14091 (W12694, W14373);
not G14092 (W12695, W14374);
not G14093 (W12696, W14375);
not G14094 (W12697, W14376);
not G14095 (W12698, W14377);
not G14096 (W12699, W14378);
not G14097 (W12700, W14379);
not G14098 (W12701, W14380);
not G14099 (W12702, W14381);
nor G14100 (W12703, W9790, W9794);
not G14101 (W12704, W14382);
not G14102 (W12705, W14383);
not G14103 (W12706, W14384);
nor G14104 (W12707, W14385, W14386);
not G14105 (W12708, W12710);
nor G14106 (W12709, W14387, W14388);
not G14107 (W12710, W14389);
nor G14108 (W12711, W14385, W14386);
not G14109 (W12712, W12714);
nor G14110 (W12713, W14390, W14391);
not G14111 (W12714, W14392);
nor G14112 (W12715, W14393, W14386);
not G14113 (W12716, W12718);
nor G14114 (W12717, W14394, W14395);
not G14115 (W12718, W14396);
nor G14116 (W12719, W14393, W14386);
not G14117 (W12720, W12722);
nor G14118 (W12721, W14397, W14398);
not G14119 (W12722, W14399);
nor G14120 (W12723, W14400, W14386);
not G14121 (W12724, W12726);
nor G14122 (W12725, W14401, W14402);
not G14123 (W12726, W14403);
nor G14124 (W12727, W11815, W12729);
and G14125 (W12728, W14404, W14405, W14406);
not G14126 (W12729, W10247);
nand G14127 (W12730, W14407, W14408);
nand G14128 (W12731, W14409, W14410);
nor G14129 (W12732, W14411, W14386);
not G14130 (W12733, W12735);
nor G14131 (W12734, W14412, W14413);
not G14132 (W12735, W14414);
nor G14133 (W12736, W14415, W14386);
not G14134 (W12737, W12739);
nor G14135 (W12738, W14416, W14417);
not G14136 (W12739, W14418);
nor G14137 (W12740, W14415, W14386);
not G14138 (W12741, W12743);
nor G14139 (W12742, W14419, W14420);
not G14140 (W12743, W14421);
not G14141 (W12744, I1005);
not G14142 (W12745, W14422);
not G14143 (W12746, W14423);
not G14144 (W12747, W14424);
nor G14145 (W12748, W14425, W14426, W14427);
not G14146 (W12749, W14428);
not G14147 (W12750, W14429);
not G14148 (W12751, W14430);
not G14149 (W12752, W8287);
not G14150 (W12753, W14431);
not G14151 (W12754, W14432);
not G14152 (W12755, W14433);
not G14153 (W12756, W11814);
not G14154 (W12757, W14434);
not G14155 (W12758, W14435);
not G14156 (W12759, W14436);
not G14157 (W12760, W14437);
not G14158 (W12761, W14438);
not G14159 (W12762, W14439);
not G14160 (W12763, W14440);
not G14161 (W12764, W14441);
not G14162 (W12765, W14442);
not G14163 (W12766, W14443);
not G14164 (W12767, W14444);
not G14165 (W12768, W14445);
not G14166 (W12769, W14446);
not G14167 (W12770, W14447);
not G14168 (W12771, W14448);
not G14169 (W12772, W14449);
not G14170 (W12773, W14450);
not G14171 (W12774, W14451);
not G14172 (W12775, W14452);
not G14173 (W12776, W14453);
not G14174 (W12777, W14454);
not G14175 (W12778, W14455);
not G14176 (W12779, W14456);
not G14177 (W12780, W14457);
not G14178 (W12781, W14458);
not G14179 (W12782, W14459);
not G14180 (W12783, W14460);
not G14181 (W12784, W14461);
not G14182 (W12785, W14462);
not G14183 (W12786, W14463);
not G14184 (W12787, W14464);
not G14185 (W12788, W14465);
not G14186 (W12789, W14466);
not G14187 (W12790, W12792);
not G14188 (W12791, I332);
not G14189 (W12792, W14467);
not G14190 (W12793, I100);
not G14191 (W12794, I333);
not G14192 (W12795, W12796);
not G14193 (W12796, W14468);
not G14194 (W12797, W12799);
not G14195 (W12798, I334);
not G14196 (W12799, W14469);
not G14197 (W12800, I335);
not G14198 (W12801, W12802);
not G14199 (W12802, W14470);
not G14200 (W12803, W12805);
not G14201 (W12804, I336);
not G14202 (W12805, W14471);
not G14203 (W12806, I337);
not G14204 (W12807, W12808);
not G14205 (W12808, W14472);
not G14206 (W12809, W12811);
not G14207 (W12810, I338);
not G14208 (W12811, W14473);
not G14209 (W12812, I339);
not G14210 (W12813, W12814);
not G14211 (W12814, W14474);
not G14212 (W12815, W12817);
not G14213 (W12816, I340);
not G14214 (W12817, W14475);
not G14215 (W12818, I341);
not G14216 (W12819, W12820);
not G14217 (W12820, W14476);
not G14218 (W12821, W13641);
and G14219 (W12822, I102, W14477);
and G14220 (W12823, W14478, W14479);
not G14221 (W12824, W14480);
and G14222 (W12825, I1423, W14481);
and G14223 (W12826, W14482, W14483);
not G14224 (W12827, W14480);
and G14225 (W12828, I1424, W14484);
and G14226 (W12829, W14485, W14486);
not G14227 (W12830, W14480);
and G14228 (W12831, I1425, W14487);
and G14229 (W12832, W14488, W14489);
not G14230 (W12833, W14480);
and G14231 (W12834, I1426, W14490);
and G14232 (W12835, W14491, W14492);
not G14233 (W12836, W14480);
not G14234 (W12837, W14493);
not G14235 (W12838, W10244);
not G14236 (W12839, W10242);
not G14237 (W12840, W10243);
not G14238 (W12841, W14494);
not G14239 (W12842, W13905);
not G14240 (W12843, W13906);
not G14241 (W12844, W13907);
not G14242 (W12845, W14495);
not G14243 (W12846, W13905);
not G14244 (W12847, W13906);
not G14245 (W12848, W13907);
and G14246 (W12849, I1427, W14496);
and G14247 (W12850, W13253, W14497);
not G14248 (W12851, I221);
not G14249 (W12852, W14498);
not G14250 (W12853, W13905);
not G14251 (W12854, W13906);
not G14252 (W12855, W13907);
not G14253 (W12856, W14499);
not G14254 (W12857, W14500);
not G14255 (W12858, W14501);
not G14256 (W12859, W14502);
and G14257 (W12860, W10243, W10207);
and G14258 (W12861, W10244, W10204);
and G14259 (W12862, W10242, W10200);
not G14260 (W12863, W5110);
not G14261 (W12864, W14500);
not G14262 (W12865, W14501);
not G14263 (W12866, W14502);
and G14264 (W12867, W10243, W10218);
and G14265 (W12868, W10244, W10215);
and G14266 (W12869, W10242, W10211);
not G14267 (W12870, W14503);
not G14268 (W12871, W14500);
not G14269 (W12872, W14501);
not G14270 (W12873, W14502);
not G14271 (W12874, W14504);
not G14272 (W12875, W14500);
not G14273 (W12876, W14501);
not G14274 (W12877, W14502);
and G14275 (W12878, W10243, W10239);
and G14276 (W12879, W10244, W10236);
and G14277 (W12880, W10242, W10232);
not G14278 (W12881, W14505);
not G14279 (W12882, W14500);
not G14280 (W12883, W14501);
not G14281 (W12884, W14502);
not G14282 (W12885, I119);
not G14283 (W12886, I118);
not G14284 (W12887, I1428);
not G14285 (W12888, W10244);
not G14286 (W12889, W10244);
and G14287 (W12890, W14506, W14507);
and G14288 (W12891, W14508, W14509);
not G14289 (W12892, W14510);
and G14290 (W12893, W14511, W14512);
and G14291 (W12894, W14513, W14514);
not G14292 (W12895, W14510);
and G14293 (W12896, I1429, W14515);
and G14294 (W12897, W14516, W14517);
not G14295 (W12898, W14510);
and G14296 (W12899, I1430, W14518);
and G14297 (W12900, W14519, W14520);
not G14298 (W12901, W14510);
and G14299 (W12902, I1431, W14521);
and G14300 (W12903, W14522, W14523);
not G14301 (W12904, W14510);
and G14302 (W12905, I1432, W14524);
and G14303 (W12906, W14525, W14526);
not G14304 (W12907, W14510);
and G14305 (W12908, I1040, W14527);
and G14306 (W12909, W14528, W14529);
not G14307 (W12910, W14530);
not G14308 (W12911, W14531);
not G14309 (W12912, W14532);
not G14310 (W12913, W14533);
not G14311 (W12914, W14534);
nor G14312 (W12915, W14535, W14536);
not G14313 (W12916, W14537);
not G14314 (W12917, W14538);
not G14315 (W12918, W10653);
nor G14316 (W12919, W14539, W14540);
not G14317 (W12920, W14537);
not G14318 (W12921, W14538);
not G14319 (W12922, W10653);
nor G14320 (W12923, W14541, W14542);
not G14321 (W12924, W14537);
not G14322 (W12925, W14538);
not G14323 (W12926, W10653);
nor G14324 (W12927, W14543, W14544);
not G14325 (W12928, W14537);
not G14326 (W12929, W14538);
not G14327 (W12930, W10653);
nor G14328 (W12931, W14545, W14546);
not G14329 (W12932, W14537);
not G14330 (W12933, W14538);
not G14331 (W12934, W10653);
nor G14332 (W12935, W14547, W14548);
not G14333 (W12936, W14537);
not G14334 (W12937, W14538);
not G14335 (W12938, W10653);
nor G14336 (W12939, W14549, W14550);
not G14337 (W12940, W10653);
not G14338 (W12941, W14537);
not G14339 (W12942, W14538);
nor G14340 (W12943, W14551, W14552);
not G14341 (W12944, W10653);
not G14342 (W12945, W14537);
not G14343 (W12946, W14538);
nor G14344 (W12947, W14553, W14554);
not G14345 (W12948, W14538);
not G14346 (W12949, W10653);
not G14347 (W12950, W14537);
nor G14348 (W12951, W14555, W14556);
not G14349 (W12952, W14537);
not G14350 (W12953, W14538);
not G14351 (W12954, W10653);
nor G14352 (W12955, W14557, W14558);
not G14353 (W12956, W13022);
not G14354 (W12957, W13023);
not G14355 (W12958, W13024);
nor G14356 (W12959, W14557, W14559);
not G14357 (W12960, W13022);
not G14358 (W12961, W13023);
not G14359 (W12962, W13024);
nor G14360 (W12963, W14557, W14560);
not G14361 (W12964, W13022);
not G14362 (W12965, W13023);
not G14363 (W12966, W13024);
nor G14364 (W12967, W14561, W14562);
not G14365 (W12968, W14563);
not G14366 (W12969, W14564);
not G14367 (W12970, W14565);
not G14368 (W12971, W14566);
nand G14369 (W12972, W14567, W14568);
nor G14370 (W12973, W14569, W14570, W14571);
and G14371 (W12974, W14572, W13986);
nor G14372 (W12975, W14573, W14574, W14575);
nor G14373 (W12976, W14576, W14577);
not G14374 (W12977, W14578);
or G14375 (W12978, W5115, W14579);
or G14376 (W12979, W14580, W14581, W5123);
or G14377 (W12980, W14582, W14581, W14583);
not G14378 (W12981, W14584);
nor G14379 (W12982, W14585, W14586);
nor G14380 (W12983, W14587, W14588);
not G14381 (W12984, W14589);
or G14382 (W12985, W14590, W14582, W5123);
or G14383 (W12986, W14590, W14580, W14583);
not G14384 (W12987, W14591);
not G14385 (W12988, W14592);
not G14386 (W12989, W14593);
not G14387 (W12990, W14594);
not G14388 (W12991, W14595);
not G14389 (W12992, W14596);
not G14390 (W12993, W14597);
not G14391 (W12994, W14598);
not G14392 (W12995, W14599);
nand G14393 (W12996, W14600, W14601);
not G14394 (W12997, W13022);
not G14395 (W12998, W13023);
not G14396 (W12999, W13024);
not G14397 (W13000, I1433);
not G14398 (W13001, W14602);
nor G14399 (W13002, W14603, W14604);
not G14400 (W13003, W14605);
not G14401 (W13004, W14606);
not G14402 (W13005, W14607);
not G14403 (W13006, W14608);
not G14404 (W13007, W13024);
not G14405 (W13008, W13022);
not G14406 (W13009, W13023);
nand G14407 (W13010, W14609, W14610);
not G14408 (W13011, W13022);
not G14409 (W13012, W13023);
not G14410 (W13013, W13024);
nand G14411 (W13014, W14611, W14612);
not G14412 (W13015, W13022);
not G14413 (W13016, W13023);
not G14414 (W13017, W13024);
not G14415 (W13018, W14613);
not G14416 (W13019, W14614);
not G14417 (W13020, W14615);
not G14418 (W13021, W14616);
not G14419 (W13022, W14617);
not G14420 (W13023, W14618);
not G14421 (W13024, W14619);
not G14422 (W13025, I242);
not G14423 (W13026, W14620);
not G14424 (W13027, I243);
not G14425 (W13028, W14621);
not G14426 (W13029, I244);
not G14427 (W13030, W14622);
not G14428 (W13031, I245);
not G14429 (W13032, W14623);
not G14430 (W13033, I246);
not G14431 (W13034, W14624);
nor G14432 (W13035, W14625, W14626, W14627);
not G14433 (W13036, W14628);
not G14434 (W13037, I239);
not G14435 (W13038, W14629);
nor G14436 (W13039, W14630, W14631, W14632);
not G14437 (W13040, W14633);
not G14438 (W13041, I240);
not G14439 (W13042, W14634);
not G14440 (W13043, I241);
not G14441 (W13044, W14635);
not G14442 (W13045, W14636);
not G14443 (W13046, W14637);
not G14444 (W13047, W14638);
not G14445 (W13048, W14639);
not G14446 (W13049, W14640);
not G14447 (W13050, W14641);
not G14448 (W13051, W14642);
not G14449 (W13052, W14643);
not G14450 (W13053, W14644);
not G14451 (W13054, W14645);
not G14452 (W13055, W14646);
not G14453 (W13056, W14647);
not G14454 (W13057, W14648);
not G14455 (W13058, W14649);
not G14456 (W13059, W14650);
not G14457 (W13060, W14651);
not G14458 (W13061, W14652);
not G14459 (W13062, W14653);
not G14460 (W13063, W14654);
not G14461 (W13064, W14655);
not G14462 (W13065, W13067);
not G14463 (W13066, I1142);
not G14464 (W13067, W14656);
not G14465 (W13068, I1434);
not G14466 (W13069, I1435);
not G14467 (W13070, W13986);
not G14468 (W13071, I1143);
not G14469 (W13072, W13073);
not G14470 (W13073, W14657);
not G14471 (W13074, W13076);
not G14472 (W13075, I1144);
not G14473 (W13076, W14658);
not G14474 (W13077, I1145);
not G14475 (W13078, W13079);
not G14476 (W13079, W14659);
not G14477 (W13080, W13082);
not G14478 (W13081, I1146);
not G14479 (W13082, W14660);
not G14480 (W13083, I1147);
not G14481 (W13084, W13085);
not G14482 (W13085, W14661);
not G14483 (W13086, W13088);
not G14484 (W13087, I1148);
not G14485 (W13088, W14662);
not G14486 (W13089, I1149);
not G14487 (W13090, W13091);
not G14488 (W13091, W14663);
not G14489 (W13092, W13094);
not G14490 (W13093, I1150);
not G14491 (W13094, W14664);
not G14492 (W13095, I1151);
not G14493 (W13096, W13097);
not G14494 (W13097, W14665);
and G14495 (W13098, W10575, W10583, W10587, W10551);
and G14496 (W13099, W10555, W10559, W10563, W10567);
not G14497 (W13100, W14666);
not G14498 (W13101, W14667);
not G14499 (W13102, W14668);
not G14500 (W13103, W14669);
not G14501 (W13104, W14670);
not G14502 (W13105, W14671);
not G14503 (W13106, W14672);
not G14504 (W13107, W14673);
not G14505 (W13108, W14674);
nor G14506 (W13109, W10559, W10563);
not G14507 (W13110, W14675);
not G14508 (W13111, W14676);
not G14509 (W13112, W14677);
nor G14510 (W13113, W14678, W14679);
not G14511 (W13114, W13116);
nor G14512 (W13115, W14680, W14681);
not G14513 (W13116, W14682);
nor G14514 (W13117, W14678, W14679);
not G14515 (W13118, W13120);
nor G14516 (W13119, W14683, W14684);
not G14517 (W13120, W14685);
nor G14518 (W13121, W14686, W14679);
not G14519 (W13122, W13124);
nor G14520 (W13123, W14687, W14688);
not G14521 (W13124, W14689);
nor G14522 (W13125, W14686, W14679);
not G14523 (W13126, W13128);
nor G14524 (W13127, W14690, W14691);
not G14525 (W13128, W14692);
nor G14526 (W13129, W14693, W14679);
not G14527 (W13130, W13132);
nor G14528 (W13131, W14694, W14695);
not G14529 (W13132, W14696);
nor G14530 (W13133, W11788, W13135);
and G14531 (W13134, W14697, W14698, W14699);
not G14532 (W13135, W11020);
nand G14533 (W13136, W14700, W14701);
nand G14534 (W13137, W14702, W14703);
nor G14535 (W13138, W14704, W14679);
not G14536 (W13139, W13141);
nor G14537 (W13140, W14705, W14706);
not G14538 (W13141, W14707);
nor G14539 (W13142, W14708, W14679);
not G14540 (W13143, W13145);
nor G14541 (W13144, W14709, W14710);
not G14542 (W13145, W14711);
nor G14543 (W13146, W14708, W14679);
not G14544 (W13147, W13149);
nor G14545 (W13148, W14712, W14713);
not G14546 (W13149, W14714);
not G14547 (W13150, I1206);
not G14548 (W13151, W14715);
not G14549 (W13152, W14716);
not G14550 (W13153, W14717);
nor G14551 (W13154, W14718, W14719, W14720);
not G14552 (W13155, W14721);
not G14553 (W13156, W14722);
not G14554 (W13157, W14723);
not G14555 (W13158, W8244);
not G14556 (W13159, W14724);
not G14557 (W13160, W14725);
not G14558 (W13161, W14726);
not G14559 (W13162, W11787);
not G14560 (W13163, W14727);
not G14561 (W13164, W14728);
not G14562 (W13165, W14729);
not G14563 (W13166, W14730);
not G14564 (W13167, W14731);
not G14565 (W13168, W14732);
not G14566 (W13169, W14733);
not G14567 (W13170, W14734);
not G14568 (W13171, W14735);
not G14569 (W13172, W14736);
not G14570 (W13173, W14737);
not G14571 (W13174, W14738);
not G14572 (W13175, W14739);
not G14573 (W13176, W14740);
not G14574 (W13177, W14741);
not G14575 (W13178, W14742);
not G14576 (W13179, W14743);
not G14577 (W13180, W14744);
not G14578 (W13181, W14745);
not G14579 (W13182, W14746);
not G14580 (W13183, W14747);
not G14581 (W13184, W14748);
not G14582 (W13185, W14749);
not G14583 (W13186, W14750);
not G14584 (W13187, W14751);
not G14585 (W13188, W14752);
not G14586 (W13189, W14753);
not G14587 (W13190, W14754);
not G14588 (W13191, W14755);
not G14589 (W13192, W14756);
not G14590 (W13193, W14757);
not G14591 (W13194, W14758);
not G14592 (W13195, W14759);
not G14593 (W13196, W13198);
not G14594 (W13197, I368);
not G14595 (W13198, W14760);
not G14596 (W13199, I149);
not G14597 (W13200, I369);
not G14598 (W13201, W13202);
not G14599 (W13202, W14761);
not G14600 (W13203, W13205);
not G14601 (W13204, I370);
not G14602 (W13205, W14762);
not G14603 (W13206, I371);
not G14604 (W13207, W13208);
not G14605 (W13208, W14763);
not G14606 (W13209, W13211);
not G14607 (W13210, I372);
not G14608 (W13211, W14764);
not G14609 (W13212, I373);
not G14610 (W13213, W13214);
not G14611 (W13214, W14765);
not G14612 (W13215, W13217);
not G14613 (W13216, I374);
not G14614 (W13217, W14766);
not G14615 (W13218, I375);
not G14616 (W13219, W13220);
not G14617 (W13220, W14767);
not G14618 (W13221, W13223);
not G14619 (W13222, I376);
not G14620 (W13223, W14768);
not G14621 (W13224, I377);
not G14622 (W13225, W13226);
not G14623 (W13226, W14769);
not G14624 (W13227, W13640);
and G14625 (W13228, I151, W14770);
not G14626 (W13229, W14771);
not G14627 (W13230, W14772);
and G14628 (W13231, I1436, W14773);
not G14629 (W13232, W14772);
and G14630 (W13233, I1437, W14774);
not G14631 (W13234, W14772);
and G14632 (W13235, I1438, W14775);
not G14633 (W13236, W14772);
and G14634 (W13237, I1439, W14776);
not G14635 (W13238, W14772);
not G14636 (W13239, W14777);
not G14637 (W13240, W11017);
not G14638 (W13241, W11015);
not G14639 (W13242, W11016);
not G14640 (W13243, W14778);
not G14641 (W13244, W13905);
not G14642 (W13245, W13906);
not G14643 (W13246, W13907);
not G14644 (W13247, W14779);
not G14645 (W13248, W13905);
not G14646 (W13249, W13906);
not G14647 (W13250, W13907);
and G14648 (W13251, I1440, W14780);
not G14649 (W13252, I222);
not G14650 (W13253, W14781);
not G14651 (W13254, W13905);
not G14652 (W13255, W13906);
not G14653 (W13256, W13907);
not G14654 (W13257, W14782);
not G14655 (W13258, W14783);
not G14656 (W13259, W14784);
not G14657 (W13260, W14785);
and G14658 (W13261, W11016, W10980);
and G14659 (W13262, W11017, W10977);
and G14660 (W13263, W11015, W10973);
not G14661 (W13264, W5385);
not G14662 (W13265, W14783);
not G14663 (W13266, W14784);
not G14664 (W13267, W14785);
and G14665 (W13268, W11016, W10991);
and G14666 (W13269, W11017, W10988);
and G14667 (W13270, W11015, W10984);
not G14668 (W13271, W14786);
not G14669 (W13272, W14783);
not G14670 (W13273, W14784);
not G14671 (W13274, W14785);
not G14672 (W13275, W14787);
not G14673 (W13276, W14783);
not G14674 (W13277, W14784);
not G14675 (W13278, W14785);
and G14676 (W13279, W11016, W11012);
and G14677 (W13280, W11017, W11009);
and G14678 (W13281, W11015, W11005);
not G14679 (W13282, W14788);
not G14680 (W13283, W14783);
not G14681 (W13284, W14784);
not G14682 (W13285, W14785);
not G14683 (W13286, I168);
not G14684 (W13287, I167);
not G14685 (W13288, I1441);
not G14686 (W13289, W11017);
not G14687 (W13290, W11017);
and G14688 (W13291, W14789, W14790);
not G14689 (W13292, W14791);
and G14690 (W13293, W14792, W14793);
not G14691 (W13294, W14791);
and G14692 (W13295, I1442, W14794);
not G14693 (W13296, W14791);
and G14694 (W13297, I1443, W14795);
not G14695 (W13298, W14791);
and G14696 (W13299, I1444, W14796);
not G14697 (W13300, W14791);
and G14698 (W13301, I1445, W14797);
not G14699 (W13302, W14791);
and G14700 (W13303, I1241, W14798);
and G14701 (W13304, W14799, W14800);
not G14702 (W13305, W14801);
not G14703 (W13306, W14802);
not G14704 (W13307, W14803);
not G14705 (W13308, W14804);
not G14706 (W13309, W14805);
nor G14707 (W13310, W14806, W14807);
not G14708 (W13311, W14808);
not G14709 (W13312, W14809);
not G14710 (W13313, W11426);
nor G14711 (W13314, W14810, W14811);
not G14712 (W13315, W14808);
not G14713 (W13316, W14809);
not G14714 (W13317, W11426);
nor G14715 (W13318, W14812, W14813);
not G14716 (W13319, W14808);
not G14717 (W13320, W14809);
not G14718 (W13321, W11426);
nor G14719 (W13322, W14814, W14815);
not G14720 (W13323, W14808);
not G14721 (W13324, W14809);
not G14722 (W13325, W11426);
nor G14723 (W13326, W14816, W14817);
not G14724 (W13327, W14808);
not G14725 (W13328, W14809);
not G14726 (W13329, W11426);
nor G14727 (W13330, W14818, W14819);
not G14728 (W13331, W14808);
not G14729 (W13332, W14809);
not G14730 (W13333, W11426);
nor G14731 (W13334, W14820, W14821);
not G14732 (W13335, W14808);
not G14733 (W13336, W14809);
not G14734 (W13337, W11426);
nor G14735 (W13338, W14822, W14823);
not G14736 (W13339, W14808);
not G14737 (W13340, W14809);
not G14738 (W13341, W11426);
nor G14739 (W13342, W14824, W14825);
not G14740 (W13343, W11426);
not G14741 (W13344, W14808);
not G14742 (W13345, W14809);
nor G14743 (W13346, W14826, W14827);
not G14744 (W13347, W14809);
not G14745 (W13348, W11426);
not G14746 (W13349, W14808);
nor G14747 (W13350, W14828, W14829);
not G14748 (W13351, W13417);
not G14749 (W13352, W13418);
not G14750 (W13353, W13419);
nor G14751 (W13354, W14828, W14830);
not G14752 (W13355, W13417);
not G14753 (W13356, W13418);
not G14754 (W13357, W13419);
nor G14755 (W13358, W14828, W14831);
not G14756 (W13359, W13417);
not G14757 (W13360, W13418);
not G14758 (W13361, W13419);
nor G14759 (W13362, W14832, W14833);
not G14760 (W13363, W14834);
not G14761 (W13364, W14835);
not G14762 (W13365, W14836);
not G14763 (W13366, W14837);
nand G14764 (W13367, W14838, W14839);
nor G14765 (W13368, W14840, W14841, W14842);
and G14766 (W13369, W14843, W13986);
nor G14767 (W13370, W14844, W14845, W14846);
nor G14768 (W13371, W14847, W14848);
not G14769 (W13372, W14849);
or G14770 (W13373, W5390, W14850);
or G14771 (W13374, W14851, W14852, W5398);
or G14772 (W13375, W14853, W14852, W14854);
not G14773 (W13376, W14855);
nor G14774 (W13377, W14856, W14857);
nor G14775 (W13378, W14858, W14859);
not G14776 (W13379, W14860);
or G14777 (W13380, W14861, W14853, W5398);
or G14778 (W13381, W14861, W14851, W14854);
not G14779 (W13382, W14862);
not G14780 (W13383, W14863);
not G14781 (W13384, W14864);
not G14782 (W13385, W14865);
not G14783 (W13386, W14866);
not G14784 (W13387, W14867);
not G14785 (W13388, W14868);
not G14786 (W13389, W14869);
not G14787 (W13390, W14870);
nand G14788 (W13391, W14871, W14872);
not G14789 (W13392, W13417);
not G14790 (W13393, W13418);
not G14791 (W13394, W13419);
not G14792 (W13395, I1446);
not G14793 (W13396, W14873);
nor G14794 (W13397, W14874, W14875);
not G14795 (W13398, W14876);
not G14796 (W13399, W14877);
not G14797 (W13400, W14878);
not G14798 (W13401, W14879);
not G14799 (W13402, W13419);
not G14800 (W13403, W13417);
not G14801 (W13404, W13418);
nand G14802 (W13405, W14880, W14881);
not G14803 (W13406, W13417);
not G14804 (W13407, W13418);
not G14805 (W13408, W13419);
nand G14806 (W13409, W14882, W14883);
not G14807 (W13410, W13417);
not G14808 (W13411, W13418);
not G14809 (W13412, W13419);
not G14810 (W13413, W14884);
not G14811 (W13414, W14885);
not G14812 (W13415, W14886);
not G14813 (W13416, W14887);
not G14814 (W13417, W14888);
not G14815 (W13418, W14889);
not G14816 (W13419, W14890);
not G14817 (W13420, I235);
not G14818 (W13421, W14891);
not G14819 (W13422, I236);
not G14820 (W13423, W14892);
not G14821 (W13424, I237);
not G14822 (W13425, W14893);
not G14823 (W13426, I238);
not G14824 (W13427, W14894);
nor G14825 (W13428, W14895, W14896, W14897);
not G14826 (W13429, W14898);
not G14827 (W13430, I231);
not G14828 (W13431, W14899);
nor G14829 (W13432, W14900, W14901, W14902);
not G14830 (W13433, W14903);
not G14831 (W13434, I232);
not G14832 (W13435, W14904);
not G14833 (W13436, I233);
not G14834 (W13437, W14905);
not G14835 (W13438, W14906);
not G14836 (W13439, I234);
not G14837 (W13440, W14907);
not G14838 (W13441, W14908);
not G14839 (W13442, W14909);
not G14840 (W13443, W14910);
not G14841 (W13444, W14911);
not G14842 (W13445, W14912);
not G14843 (W13446, W14913);
not G14844 (W13447, W14914);
not G14845 (W13448, W14915);
not G14846 (W13449, W14916);
not G14847 (W13450, W14917);
not G14848 (W13451, W14918);
not G14849 (W13452, W14919);
not G14850 (W13453, W14920);
not G14851 (W13454, W14921);
not G14852 (W13455, W14922);
not G14853 (W13456, W14923);
not G14854 (W13457, W14924);
not G14855 (W13458, W14925);
not G14856 (W13459, W14926);
not G14857 (W13460, W13462);
not G14858 (W13461, I1343);
not G14859 (W13462, W14927);
not G14860 (W13463, I1447);
not G14861 (W13464, I1448);
not G14862 (W13465, W13986);
not G14863 (W13466, I1344);
not G14864 (W13467, W13468);
not G14865 (W13468, W14928);
not G14866 (W13469, W13471);
not G14867 (W13470, I1345);
not G14868 (W13471, W14929);
not G14869 (W13472, I1346);
not G14870 (W13473, W13474);
not G14871 (W13474, W14930);
not G14872 (W13475, W13477);
not G14873 (W13476, I1347);
not G14874 (W13477, W14931);
not G14875 (W13478, I1348);
not G14876 (W13479, W13480);
not G14877 (W13480, W14932);
not G14878 (W13481, W13483);
not G14879 (W13482, I1349);
not G14880 (W13483, W14933);
not G14881 (W13484, I1350);
not G14882 (W13485, W13486);
not G14883 (W13486, W14934);
not G14884 (W13487, W13489);
not G14885 (W13488, I1351);
not G14886 (W13489, W14935);
not G14887 (W13490, I1352);
not G14888 (W13491, W13492);
not G14889 (W13492, W14936);
and G14890 (W13493, W11344, W11352, W11356, W11363);
and G14891 (W13494, W11324, W11328, W11332, W11336);
not G14892 (W13495, W14937);
not G14893 (W13496, W14938);
not G14894 (W13497, W14939);
not G14895 (W13498, W14940);
not G14896 (W13499, W14941);
not G14897 (W13500, W14942);
not G14898 (W13501, W14943);
not G14899 (W13502, W14944);
not G14900 (W13503, W14945);
nor G14901 (W13504, W11328, W11332);
not G14902 (W13505, W14946);
not G14903 (W13506, W14947);
not G14904 (W13507, W14948);
not G14905 (W13508, W14949);
not G14906 (W13509, W14950);
nand G14907 (W13510, W11616, W14951);
nand G14908 (W13511, W14952, W14951);
not G14909 (W13512, W14953);
not G14910 (W13513, W14954);
nand G14911 (W13514, W11618, W14955);
nand G14912 (W13515, W14952, W14955);
not G14913 (W13516, W14954);
not G14914 (W13517, W14953);
not G14915 (W13518, W14956);
not G14916 (W13519, W14957);
not G14917 (W13520, W14958);
not G14918 (W13521, W14959);
not G14919 (W13522, W14954);
not G14920 (W13523, W14954);
not G14921 (W13524, W14954);
not G14922 (W13525, W14954);
not G14923 (W13526, W14954);
not G14924 (W13527, W14954);
not G14925 (W13528, W14954);
not G14926 (W13529, W14954);
not G14927 (W13530, W14953);
not G14928 (W13531, W14953);
not G14929 (W13532, W14953);
not G14930 (W13533, W14953);
not G14931 (W13534, W14953);
not G14932 (W13535, W14953);
not G14933 (W13536, W14953);
not G14934 (W13537, W14953);
not G14935 (W13538, W14953);
not G14936 (W13539, W14953);
not G14937 (W13540, W14953);
not G14938 (W13541, W14953);
not G14939 (W13542, W14953);
not G14940 (W13543, W14953);
not G14941 (W13544, W14953);
not G14942 (W13545, W14953);
not G14943 (W13546, W14954);
not G14944 (W13547, W14954);
not G14945 (W13548, W14954);
not G14946 (W13549, W14954);
not G14947 (W13550, W14954);
not G14948 (W13551, W14954);
not G14949 (W13552, W14954);
not G14950 (W13553, W14954);
nand G14951 (W13554, W14960, W14961);
nand G14952 (W13555, W14962, W14961);
nand G14953 (W13556, W14963, W14964);
nand G14954 (W13557, W14965, W14964);
not G14955 (W13558, W14966);
not G14956 (W13559, I1381);
not G14957 (W13560, W13561);
not G14958 (W13561, W14967);
not G14959 (W13562, I1382);
not G14960 (W13563, W13564);
not G14961 (W13564, W14968);
not G14962 (W13565, W13567);
not G14963 (W13566, I1383);
not G14964 (W13567, W14969);
not G14965 (W13568, W13570);
not G14966 (W13569, I1384);
not G14967 (W13570, W14970);
and G14968 (W13571, W11644, I1384, W13562);
not G14969 (W13572, W13574);
not G14970 (W13573, I1385);
not G14971 (W13574, W14971);
not G14972 (W13575, I1386);
not G14973 (W13576, W13577);
not G14974 (W13577, W14972);
not G14975 (W13578, W13580);
not G14976 (W13579, I1387);
not G14977 (W13580, W14973);
not G14978 (W13581, I1388);
not G14979 (W13582, W13583);
not G14980 (W13583, W14974);
not G14981 (W13584, W13586);
not G14982 (W13585, I1389);
not G14983 (W13586, W14975);
not G14984 (W13587, I1390);
not G14985 (W13588, W13589);
not G14986 (W13589, W14976);
not G14987 (W13590, W13592);
not G14988 (W13591, I1391);
not G14989 (W13592, W14977);
and G14990 (W13593, W14978, W13591, I1386, W13579);
and G14991 (W13594, I1388, I1389, W13587, I1385);
not G14992 (W13595, W14979);
not G14993 (W13596, I412);
not G14994 (W13597, W14980);
not G14995 (W13598, W14981);
nand G14996 (W13599, W14982, W14983);
nand G14997 (W13600, W13599, W13601);
nand G14998 (W13601, W14984, W14985);
not G14999 (W13602, W14986);
nand G15000 (W13603, W14987, W14988);
nand G15001 (W13604, W13603, W13605);
nand G15002 (W13605, W14989, W14990);
not G15003 (W13606, W14991);
not G15004 (W13607, W14992);
and G15005 (W13608, W14993, W14994);
and G15006 (W13609, W14995, W14996);
and G15007 (W13610, W14997, W14998);
and G15008 (W13611, W14999, W15000);
not G15009 (W13612, W15001);
nor G15010 (W13613, W15002, W15003);
nor G15011 (W13614, W15004, W15005);
and G15012 (W13615, W15006, W15007);
and G15013 (W13616, W15008, W15009);
and G15014 (W13617, W15010, W15011);
and G15015 (W13618, W15012, W15013);
not G15016 (W13619, W15014);
nor G15017 (W13620, W15015, W15016);
nor G15018 (W13621, W15017, W15018);
and G15019 (W13622, W15019, W15020);
and G15020 (W13623, W15021, W15022);
and G15021 (W13624, W15023, W15024);
and G15022 (W13625, W15025, W15026);
not G15023 (W13626, W15027);
nor G15024 (W13627, W15028, W15029);
nor G15025 (W13628, W15030, W15031);
and G15026 (W13629, W15032, W15033);
and G15027 (W13630, W15034, W15035);
and G15028 (W13631, W15036, W15037);
and G15029 (W13632, W15038, W15039);
not G15030 (W13633, W15040);
nor G15031 (W13634, W15041, W15042);
nor G15032 (W13635, W15043, W15044);
not G15033 (W13636, W15045);
not G15034 (W13637, W15046);
not G15035 (W13638, W15047);
not G15036 (W13639, W11874);
not G15037 (W13640, W15048);
not G15038 (W13641, W15049);
not G15039 (W13642, W15050);
not G15040 (W13643, W15051);
and G15041 (W13644, W13651, W5250);
and G15042 (W13645, W13653, W15052, W5253);
and G15043 (W13646, W13653, W13652, W5252);
and G15044 (W13647, W15053, W5251);
and G15045 (W13648, W15053, W15052, W13650);
nand G15046 (W13649, W15054, W11017);
not G15047 (W13650, W5252);
not G15048 (W13651, W13653);
not G15049 (W13652, W5251);
not G15050 (W13653, W15055);
not G15051 (W13654, W5253);
nand G15052 (W13655, W15054, W11017);
and G15053 (W13656, W13651, W5252, W13654);
and G15054 (W13657, W13653, W5252, W5253);
and G15055 (W13658, W15056, W13653, W13654);
and G15056 (W13659, W15056, W13651, W5253);
nand G15057 (W13660, W15054, W11017);
nand G15058 (W13661, W13650, W13652);
nand G15059 (W13662, W15054, W11017);
nand G15060 (W13663, W15054, W11016);
nand G15061 (W13664, W15054, W11015);
nand G15062 (W13665, W15054, W11016);
nand G15063 (W13666, W15054, W11015);
nand G15064 (W13667, W15054, W11016);
nand G15065 (W13668, W15054, W11015);
nand G15066 (W13669, W15054, W11016);
nand G15067 (W13670, W15054, W11015);
nor G15068 (W13671, W15057, W15058, W15059);
and G15069 (W13672, W11890, W11872, W15060);
and G15070 (W13673, W11015, I1214);
and G15071 (W13674, W11016, I1215);
and G15072 (W13675, W11017, I1213);
and G15073 (W13676, W11015, I452);
and G15074 (W13677, W11016, I453);
and G15075 (W13678, W11017, I454);
and G15076 (W13679, W13686, W4975);
and G15077 (W13680, W13688, W15061, W4978);
and G15078 (W13681, W13688, W13687, W4977);
and G15079 (W13682, W15062, W4976);
and G15080 (W13683, W15062, W15061, W13685);
nand G15081 (W13684, W15063, W10244);
not G15082 (W13685, W4977);
not G15083 (W13686, W13688);
not G15084 (W13687, W4976);
not G15085 (W13688, W15055);
not G15086 (W13689, W4978);
nand G15087 (W13690, W15063, W10244);
and G15088 (W13691, W13686, W4977, W13689);
and G15089 (W13692, W13688, W4977, W4978);
and G15090 (W13693, W15064, W13688, W13689);
and G15091 (W13694, W15064, W13686, W4978);
nand G15092 (W13695, W15063, W10244);
nand G15093 (W13696, W13685, W13687);
nand G15094 (W13697, W15063, W10244);
nand G15095 (W13698, W15063, W10243);
nand G15096 (W13699, W15063, W10242);
nand G15097 (W13700, W15063, W10243);
nand G15098 (W13701, W15063, W10242);
nand G15099 (W13702, W15063, W10243);
nand G15100 (W13703, W15063, W10242);
nand G15101 (W13704, W15063, W10243);
nand G15102 (W13705, W15063, W10242);
nor G15103 (W13706, W15065, W15066, W15067);
and G15104 (W13707, W10242, I1013);
and G15105 (W13708, W10243, I1014);
and G15106 (W13709, W10244, I1012);
and G15107 (W13710, W10242, I464);
and G15108 (W13711, W10243, I465);
and G15109 (W13712, W10244, I466);
and G15110 (W13713, W13720, W4700);
and G15111 (W13714, W13722, W15068, W4703);
and G15112 (W13715, W13722, W13721, W4702);
and G15113 (W13716, W15069, W4701);
and G15114 (W13717, W15069, W15068, W13719);
nand G15115 (W13718, W15070, W9471);
not G15116 (W13719, W4702);
not G15117 (W13720, W13722);
not G15118 (W13721, W4701);
not G15119 (W13722, W15055);
not G15120 (W13723, W4703);
nand G15121 (W13724, W15070, W9471);
and G15122 (W13725, W13720, W4702, W13723);
and G15123 (W13726, W13722, W4702, W4703);
and G15124 (W13727, W15071, W13722, W13723);
and G15125 (W13728, W15071, W13720, W4703);
nand G15126 (W13729, W15070, W9471);
nand G15127 (W13730, W13719, W13721);
nand G15128 (W13731, W15070, W9471);
nand G15129 (W13732, W15070, W9470);
nand G15130 (W13733, W15070, W9469);
nand G15131 (W13734, W15070, W9470);
nand G15132 (W13735, W15070, W9469);
nand G15133 (W13736, W15070, W9470);
nand G15134 (W13737, W15070, W9469);
nand G15135 (W13738, W15070, W9470);
nand G15136 (W13739, W15070, W9469);
nor G15137 (W13740, W15072, W15073, W15074);
and G15138 (W13741, W9469, I812);
and G15139 (W13742, W9470, I813);
and G15140 (W13743, W9471, I811);
and G15141 (W13744, W9469, I476);
and G15142 (W13745, W9470, I477);
and G15143 (W13746, W9471, I478);
and G15144 (W13747, W13754, W4425);
and G15145 (W13748, W13756, W15075, W4428);
and G15146 (W13749, W13756, W13755, W4427);
and G15147 (W13750, W15076, W4426);
and G15148 (W13751, W15076, W15075, W13753);
nand G15149 (W13752, W15077, W8698);
not G15150 (W13753, W4427);
not G15151 (W13754, W13756);
not G15152 (W13755, W4426);
not G15153 (W13756, W15055);
not G15154 (W13757, W4428);
nand G15155 (W13758, W15077, W8698);
and G15156 (W13759, W13754, W4427, W13757);
and G15157 (W13760, W13756, W4427, W4428);
and G15158 (W13761, W15078, W13756, W13757);
and G15159 (W13762, W15078, W13754, W4428);
nand G15160 (W13763, W15077, W8698);
nand G15161 (W13764, W13753, W13755);
nand G15162 (W13765, W15077, W8698);
nand G15163 (W13766, W15077, W8697);
nand G15164 (W13767, W15077, W8696);
nand G15165 (W13768, W15077, W8697);
nand G15166 (W13769, W15077, W8696);
nand G15167 (W13770, W15077, W8697);
nand G15168 (W13771, W15077, W8696);
nand G15169 (W13772, W15077, W8697);
nand G15170 (W13773, W15077, W8696);
nor G15171 (W13774, W15079, W15080, W15081);
and G15172 (W13775, W8696, I611);
and G15173 (W13776, W8697, I612);
and G15174 (W13777, W8698, I610);
and G15175 (W13778, W8696, I488);
and G15176 (W13779, W8697, I489);
and G15177 (W13780, W8698, I490);
not G15178 (W13781, W15082);
and G15179 (W13782, I559, W11890, I556, W15083);
not G15180 (W13783, W5846);
not G15181 (W13784, W13786);
not G15182 (W13785, I1395);
not G15183 (W13786, W15084);
not G15184 (W13787, I1396);
not G15185 (W13788, W13789);
not G15186 (W13789, W15085);
not G15187 (W13790, W15086);
not G15188 (W13791, W15087);
not G15189 (W13792, W15088);
not G15190 (W13793, W15089);
not G15191 (W13794, W15090);
nor G15192 (W13795, W15091, W15092);
not G15193 (W13796, W15093);
and G15194 (W13797, W15094, W15095);
and G15195 (W13798, W15096, W15097);
not G15196 (W13799, W13816);
and G15197 (W13800, W15098, W15099);
and G15198 (W13801, W15100, W15101);
not G15199 (W13802, W13816);
nor G15200 (W13803, W15091, W15102);
and G15201 (W13804, W15103, W15104);
and G15202 (W13805, W15105, W15106);
not G15203 (W13806, W13816);
and G15204 (W13807, W15107, W15108);
and G15205 (W13808, W15109, W15110);
not G15206 (W13809, W13816);
nor G15207 (W13810, W15111, W15091, W15112);
and G15208 (W13811, W15113, W15114);
and G15209 (W13812, W15115, W15116);
not G15210 (W13813, W13816);
nor G15211 (W13814, W15117, W15091);
not G15212 (W13815, W15118);
not G15213 (W13816, W15119);
nand G15214 (W13817, W13821, W15120);
nand G15215 (W13818, W13810, W15120);
nand G15216 (W13819, W15121, W15122);
nand G15217 (W13820, W15123, W15122);
nor G15218 (W13821, W15111, W15091, W15124);
and G15219 (W13822, W15125, W15126);
and G15220 (W13823, W15127, W15128);
not G15221 (W13824, W13816);
not G15222 (W13825, W15091);
and G15223 (W13826, W15129, W15130);
and G15224 (W13827, W15131, W15132);
not G15225 (W13828, W13816);
and G15226 (W13829, W15133, W15134);
and G15227 (W13830, W15135, W15136);
not G15228 (W13831, W13816);
nand G15229 (W13832, W15137, W13643);
nand G15230 (W13833, W15137, W8544);
nand G15231 (W13834, W15137, W15138);
not G15232 (W13835, W15139);
not G15233 (W13836, W15140);
and G15234 (W13837, W15141, W15142);
nand G15235 (W13838, W15143, W13643);
nand G15236 (W13839, W15143, W8544);
nand G15237 (W13840, W15143, W15138);
nand G15238 (W13841, W8412, W13643);
nand G15239 (W13842, W8412, W8544);
nand G15240 (W13843, W8412, W15138);
nand G15241 (W13844, W8412, W13643);
nand G15242 (W13845, W8412, W8544);
nand G15243 (W13846, W8412, W15138);
nand G15244 (W13847, W15143, W13643);
nand G15245 (W13848, W15143, W8544);
nand G15246 (W13849, W15143, W15138);
nand G15247 (W13850, W15143, W13643);
nand G15248 (W13851, W15143, W8544);
nand G15249 (W13852, W15143, W15138);
nand G15250 (W13853, W15143, W13643);
nand G15251 (W13854, W15143, W8544);
nand G15252 (W13855, W15143, W15138);
nand G15253 (W13856, W15143, W13643);
nand G15254 (W13857, W15143, W8544);
nand G15255 (W13858, W15143, W15138);
nand G15256 (W13859, W15143, W13643);
nand G15257 (W13860, W15143, W8544);
nand G15258 (W13861, W15143, W15138);
nand G15259 (W13862, W15143, W13643);
nand G15260 (W13863, W15143, W8544);
nand G15261 (W13864, W15143, W15138);
nand G15262 (W13865, W15143, W13643);
nand G15263 (W13866, W15143, W8544);
nand G15264 (W13867, W15143, W15138);
nand G15265 (W13868, W15143, W13643);
nand G15266 (W13869, W15143, W8544);
nand G15267 (W13870, W15143, W15138);
nand G15268 (W13871, W15143, W13643);
nand G15269 (W13872, W15143, W8544);
nand G15270 (W13873, W15143, W15138);
nand G15271 (W13874, W15143, W13643);
nand G15272 (W13875, W15143, W8544);
nand G15273 (W13876, W15143, W15138);
not G15274 (W13877, W15144);
not G15275 (W13878, W15145);
not G15276 (W13879, W15146);
not G15277 (W13880, W15147);
not G15278 (W13881, W15148);
not G15279 (W13882, W15149);
not G15280 (W13883, W15150);
not G15281 (W13884, W15151);
not G15282 (W13885, W15152);
not G15283 (W13886, W15153);
not G15284 (W13887, W13889);
not G15285 (W13888, W15154);
not G15286 (W13889, W15155);
not G15287 (W13890, W15156);
not G15288 (W13891, W13893);
not G15289 (W13892, W15157);
not G15290 (W13893, W15158);
not G15291 (W13894, W13896);
not G15292 (W13895, W15159);
not G15293 (W13896, W15160);
not G15294 (W13897, W13899);
not G15295 (W13898, W15161);
not G15296 (W13899, W15162);
not G15297 (W13900, W13902);
not G15298 (W13901, W15163);
not G15299 (W13902, W15164);
nand G15300 (W13903, W15165, W15166);
not G15301 (W13904, I1449);
not G15302 (W13905, W15167);
not G15303 (W13906, W15168);
not G15304 (W13907, W15169);
not G15305 (W13908, I219);
not G15306 (W13909, W13910);
not G15307 (W13910, W15170);
not G15308 (W13911, W4435);
not G15309 (W13912, W15171);
not G15310 (W13913, W15172);
not G15311 (W13914, W15173);
not G15312 (W13915, W15174);
not G15313 (W13916, W15175);
not G15314 (W13917, W12161);
not G15315 (W13918, W15176);
not G15316 (W13919, W15177);
not G15317 (W13920, W13922);
not G15318 (W13921, W15178);
not G15319 (W13922, W15179);
not G15320 (W13923, I1450);
not G15321 (W13924, W15180);
not G15322 (W13925, W13927);
not G15323 (W13926, W15181);
not G15324 (W13927, W15182);
not G15325 (W13928, W13930);
not G15326 (W13929, W15183);
not G15327 (W13930, W15184);
not G15328 (W13931, W13933);
not G15329 (W13932, W15185);
not G15330 (W13933, W15186);
not G15331 (W13934, W13936);
not G15332 (W13935, W15187);
not G15333 (W13936, W15188);
not G15334 (W13937, W13939);
not G15335 (W13938, W15189);
not G15336 (W13939, W15190);
not G15337 (W13940, W13942);
not G15338 (W13941, I1451);
not G15339 (W13942, W15191);
not G15340 (W13943, W15192);
nand G15341 (W13944, W15193, W15194, W9108);
nand G15342 (W13945, W15195, W12210);
nand G15343 (W13946, W15195, W12211);
nand G15344 (W13947, W15195, W12212);
and G15345 (W13948, W15196, W15197);
and G15346 (W13949, W15198, W15199);
not G15347 (W13950, W15200);
not G15348 (W13951, W15201);
and G15349 (W13952, W15202, W15203);
and G15350 (W13953, W15204, W15205);
and G15351 (W13954, W15206, W15207);
and G15352 (W13955, W15208, W15209);
and G15353 (W13956, W15210, W15211);
and G15354 (W13957, W15212, W15213);
and G15355 (W13958, W15214, W15215);
and G15356 (W13959, W15216, W15217);
and G15357 (W13960, W15218, W15219);
and G15358 (W13961, W15220, W15221);
and G15359 (W13962, W15222, W15223);
and G15360 (W13963, W15224, W15225);
and G15361 (W13964, W15226, W15227);
and G15362 (W13965, W15228, W15229);
and G15363 (W13966, W15230, W15231);
and G15364 (W13967, W15232, W15233);
and G15365 (W13968, W15234, W15235);
and G15366 (W13969, W15236, W15237);
and G15367 (W13970, W13943, W12099);
nand G15368 (W13971, W15238, W15239);
not G15369 (W13972, W15240);
nand G15370 (W13973, W15241, W15242);
and G15371 (W13974, W13982, W15243);
and G15372 (W13975, W13983, W15244, W12099);
not G15373 (W13976, W15245);
nand G15374 (W13977, W15246, W12212);
nand G15375 (W13978, W15246, W12211);
nand G15376 (W13979, W15246, W12210);
or G15377 (W13980, W15247, W15248);
or G15378 (W13981, W9109, W15249);
not G15379 (W13982, W15250);
not G15380 (W13983, W15251);
not G15381 (W13984, W15245);
not G15382 (W13985, W15171);
not G15383 (W13986, W15252);
and G15384 (W13987, W13994, W4561);
and G15385 (W13988, W13996, W15253, W4573);
and G15386 (W13989, W13996, W13995, W4569);
and G15387 (W13990, W15254, W4565);
and G15388 (W13991, W15254, W15253, W13993);
nand G15389 (W13992, W4529, W12212);
not G15390 (W13993, W4569);
not G15391 (W13994, W13996);
not G15392 (W13995, W4565);
not G15393 (W13996, W15055);
not G15394 (W13997, W4573);
nand G15395 (W13998, W4529, W12212);
and G15396 (W13999, W13994, W4569, W13997);
and G15397 (W14000, W13996, W4569, W4573);
and G15398 (W14001, W15255, W13996, W13997);
and G15399 (W14002, W15255, W13994, W4573);
nand G15400 (W14003, W4529, W12212);
nand G15401 (W14004, W13993, W13995);
nand G15402 (W14005, W4529, W12212);
nand G15403 (W14006, W4529, W12211);
nand G15404 (W14007, W4529, W12210);
nand G15405 (W14008, W4529, W12211);
nand G15406 (W14009, W4529, W12210);
nand G15407 (W14010, W4529, W12211);
nand G15408 (W14011, W4529, W12210);
nand G15409 (W14012, W4529, W12211);
nand G15410 (W14013, W4529, W12210);
nand G15411 (W14014, W15256, W15257);
nand G15412 (W14015, W15176, W15257);
nor G15413 (W14016, W15258, W15259, W15260);
nor G15414 (W14017, W15261, W15262, W15263);
and G15415 (W14018, W15261, W15262, W15263);
nand G15416 (W14019, W15264, W12210);
nand G15417 (W14020, W15264, W12211);
nand G15418 (W14021, W15264, W12212);
nand G15419 (W14022, W15265, W15266);
nand G15420 (W14023, W15267, W15268);
nand G15421 (W14024, W4560, W15268);
nand G15422 (W14025, W15269, W15270);
nand G15423 (W14026, W15271, W15270);
nor G15424 (W14027, W12188, W15272, W15273, W15274);
nand G15425 (W14028, W15275, W12210);
nand G15426 (W14029, W15275, W12211);
nand G15427 (W14030, W15275, W12212);
not G15428 (W14031, I46);
not G15429 (W14032, I45);
not G15430 (W14033, I1452);
nand G15431 (W14034, W15276, W9107);
nand G15432 (W14035, W15276, W9107);
nand G15433 (W14036, W15276, W9107);
nand G15434 (W14037, W15276, W9107);
nand G15435 (W14038, W15276, W9107);
nand G15436 (W14039, W15276, W9107);
and G15437 (W14040, W13950, W9145);
and G15438 (W14041, W13951, W9142);
and G15439 (W14042, W9107, W9139);
nand G15440 (W14043, W15276, W9107);
nand G15441 (W14044, W15276, W9107);
and G15442 (W14045, W13950, W9154);
and G15443 (W14046, W13951, W9151);
and G15444 (W14047, W9107, W9148);
nand G15445 (W14048, W15276, W9107);
nand G15446 (W14049, W15276, W9107);
nand G15447 (W14050, W15276, W13951);
nand G15448 (W14051, W15276, W13950);
nand G15449 (W14052, W15276, W13951);
nand G15450 (W14053, W15276, W13950);
nand G15451 (W14054, W15276, W13951);
nand G15452 (W14055, W15276, W13950);
nand G15453 (W14056, W15276, W13951);
nand G15454 (W14057, W15276, W13950);
nand G15455 (W14058, W15276, W13951);
nand G15456 (W14059, W15276, W13950);
nand G15457 (W14060, W15276, W13951);
nand G15458 (W14061, W15276, W13950);
nand G15459 (W14062, W15276, W13951);
nand G15460 (W14063, W15276, W13951);
nand G15461 (W14064, W15276, W13950);
nand G15462 (W14065, W15276, W13951);
nand G15463 (W14066, W15276, W13950);
nand G15464 (W14067, W15276, W13951);
nand G15465 (W14068, W15276, W13950);
nand G15466 (W14069, W15276, W13950);
not G15467 (W14070, W15277);
not G15468 (W14071, W15278);
not G15469 (W14072, W15279);
not G15470 (W14073, W15280);
not G15471 (W14074, W15281);
not G15472 (W14075, W15282);
not G15473 (W14076, W15283);
not G15474 (W14077, W15284);
not G15475 (W14078, W15285);
not G15476 (W14079, W15286);
nand G15477 (W14080, W15287, W9107);
nand G15478 (W14081, W15287, W13951);
nand G15479 (W14082, W15287, W13950);
nand G15480 (W14083, W15287, W9107);
nand G15481 (W14084, W15287, W13951);
nand G15482 (W14085, W15287, W13950);
nand G15483 (W14086, W15287, W9107);
nand G15484 (W14087, W15287, W13951);
nand G15485 (W14088, W15287, W13950);
nand G15486 (W14089, W15287, W9107);
nand G15487 (W14090, W15287, W13951);
nand G15488 (W14091, W15287, W13950);
nor G15489 (W14092, W15288, W15289);
not G15490 (W14093, W15290);
and G15491 (W14094, W15291, W15292);
and G15492 (W14095, W15293, W15294);
not G15493 (W14096, W14113);
and G15494 (W14097, W15295, W15296);
and G15495 (W14098, W15297, W15298);
not G15496 (W14099, W14113);
nor G15497 (W14100, W15288, W15299);
and G15498 (W14101, W15300, W15301);
and G15499 (W14102, W15302, W15303);
not G15500 (W14103, W14113);
and G15501 (W14104, W15304, W15305);
and G15502 (W14105, W15306, W15307);
not G15503 (W14106, W14113);
nor G15504 (W14107, W15308, W15288, W15309);
and G15505 (W14108, W15310, W15311);
and G15506 (W14109, W15312, W15313);
not G15507 (W14110, W14113);
nor G15508 (W14111, W15314, W15288);
not G15509 (W14112, W15315);
not G15510 (W14113, W15316);
nand G15511 (W14114, W14118, W15317);
nand G15512 (W14115, W14107, W15317);
nand G15513 (W14116, W15318, W15319);
nand G15514 (W14117, W15320, W15319);
nor G15515 (W14118, W15308, W15288, W15321);
and G15516 (W14119, W15322, W15323);
and G15517 (W14120, W15324, W15325);
not G15518 (W14121, W14113);
not G15519 (W14122, W15288);
and G15520 (W14123, W15326, W15327);
and G15521 (W14124, W15328, W15329);
not G15522 (W14125, W14113);
and G15523 (W14126, W15330, W15331);
and G15524 (W14127, W15332, W15333);
not G15525 (W14128, W14113);
nand G15526 (W14129, W15334, W13642);
nand G15527 (W14130, W15334, W9317);
nand G15528 (W14131, W15334, W15335);
not G15529 (W14132, W15336);
not G15530 (W14133, W15337);
and G15531 (W14134, W15338, W15339);
nand G15532 (W14135, W15340, W13642);
nand G15533 (W14136, W15340, W9317);
nand G15534 (W14137, W15340, W15335);
nand G15535 (W14138, W9185, W13642);
nand G15536 (W14139, W9185, W9317);
nand G15537 (W14140, W9185, W15335);
nand G15538 (W14141, W9185, W13642);
nand G15539 (W14142, W9185, W9317);
nand G15540 (W14143, W9185, W15335);
nand G15541 (W14144, W15340, W13642);
nand G15542 (W14145, W15340, W9317);
nand G15543 (W14146, W15340, W15335);
nand G15544 (W14147, W15340, W13642);
nand G15545 (W14148, W15340, W9317);
nand G15546 (W14149, W15340, W15335);
nand G15547 (W14150, W15340, W13642);
nand G15548 (W14151, W15340, W9317);
nand G15549 (W14152, W15340, W15335);
nand G15550 (W14153, W15340, W13642);
nand G15551 (W14154, W15340, W9317);
nand G15552 (W14155, W15340, W15335);
nand G15553 (W14156, W15340, W13642);
nand G15554 (W14157, W15340, W9317);
nand G15555 (W14158, W15340, W15335);
nand G15556 (W14159, W15340, W13642);
nand G15557 (W14160, W15340, W9317);
nand G15558 (W14161, W15340, W15335);
nand G15559 (W14162, W15340, W13642);
nand G15560 (W14163, W15340, W9317);
nand G15561 (W14164, W15340, W15335);
nand G15562 (W14165, W15340, W13642);
nand G15563 (W14166, W15340, W9317);
nand G15564 (W14167, W15340, W15335);
nand G15565 (W14168, W15340, W13642);
nand G15566 (W14169, W15340, W9317);
nand G15567 (W14170, W15340, W15335);
nand G15568 (W14171, W15340, W13642);
nand G15569 (W14172, W15340, W9317);
nand G15570 (W14173, W15340, W15335);
not G15571 (W14174, W15341);
not G15572 (W14175, W15342);
not G15573 (W14176, W15343);
not G15574 (W14177, W15344);
not G15575 (W14178, W15345);
not G15576 (W14179, W15346);
not G15577 (W14180, W15347);
not G15578 (W14181, W15348);
not G15579 (W14182, W15349);
not G15580 (W14183, W15350);
not G15581 (W14184, W14186);
not G15582 (W14185, W15351);
not G15583 (W14186, W15352);
not G15584 (W14187, W15353);
not G15585 (W14188, W14190);
not G15586 (W14189, W15354);
not G15587 (W14190, W15355);
not G15588 (W14191, W14193);
not G15589 (W14192, W15356);
not G15590 (W14193, W15357);
not G15591 (W14194, W14196);
not G15592 (W14195, W15358);
not G15593 (W14196, W15359);
not G15594 (W14197, W14199);
not G15595 (W14198, W15360);
not G15596 (W14199, W15361);
nand G15597 (W14200, W15362, W15363);
not G15598 (W14201, I1453);
not G15599 (W14202, I220);
not G15600 (W14203, W14204);
not G15601 (W14204, W15364);
not G15602 (W14205, W4710);
not G15603 (W14206, W15365);
not G15604 (W14207, W15366);
not G15605 (W14208, W15367);
not G15606 (W14209, W15368);
not G15607 (W14210, W15369);
not G15608 (W14211, W12567);
not G15609 (W14212, W15370);
not G15610 (W14213, W15371);
not G15611 (W14214, W14216);
not G15612 (W14215, W15372);
not G15613 (W14216, W15373);
not G15614 (W14217, I1454);
not G15615 (W14218, W15374);
not G15616 (W14219, W14221);
not G15617 (W14220, W15375);
not G15618 (W14221, W15376);
not G15619 (W14222, W14224);
not G15620 (W14223, W15377);
not G15621 (W14224, W15378);
not G15622 (W14225, W14227);
not G15623 (W14226, W15379);
not G15624 (W14227, W15380);
not G15625 (W14228, W14230);
not G15626 (W14229, W15381);
not G15627 (W14230, W15382);
not G15628 (W14231, W14233);
not G15629 (W14232, W15383);
not G15630 (W14233, W15384);
not G15631 (W14234, W14236);
not G15632 (W14235, I1455);
not G15633 (W14236, W15385);
not G15634 (W14237, W15386);
nand G15635 (W14238, W15387, W15388, W9881);
nand G15636 (W14239, W15389, W12616);
nand G15637 (W14240, W15389, W12617);
nand G15638 (W14241, W15389, W12618);
and G15639 (W14242, W15390, W15391);
and G15640 (W14243, W15392, W15393);
not G15641 (W14244, W15394);
not G15642 (W14245, W15395);
and G15643 (W14246, W15396, W15397);
and G15644 (W14247, W15398, W15399);
and G15645 (W14248, W15400, W15401);
and G15646 (W14249, W15402, W15403);
and G15647 (W14250, W15404, W15405);
and G15648 (W14251, W15406, W15407);
and G15649 (W14252, W15408, W15409);
and G15650 (W14253, W15410, W15411);
and G15651 (W14254, W15412, W15413);
and G15652 (W14255, W15414, W15415);
and G15653 (W14256, W15416, W15417);
and G15654 (W14257, W15418, W15419);
and G15655 (W14258, W15420, W15421);
and G15656 (W14259, W15422, W15423);
and G15657 (W14260, W15424, W15425);
and G15658 (W14261, W15426, W15427);
and G15659 (W14262, W15428, W15429);
and G15660 (W14263, W15430, W15431);
and G15661 (W14264, W14237, W12505);
nand G15662 (W14265, W15432, W15433);
not G15663 (W14266, W15434);
nand G15664 (W14267, W15435, W15436);
and G15665 (W14268, W14276, W15437);
and G15666 (W14269, W14277, W15438, W12505);
not G15667 (W14270, W15439);
nand G15668 (W14271, W15440, W12618);
nand G15669 (W14272, W15440, W12617);
nand G15670 (W14273, W15440, W12616);
or G15671 (W14274, W15441, W15442);
or G15672 (W14275, W9882, W15443);
not G15673 (W14276, W15444);
not G15674 (W14277, W15445);
not G15675 (W14278, W15439);
not G15676 (W14279, W15365);
and G15677 (W14280, W14287, W4836);
and G15678 (W14281, W14289, W15446, W4848);
and G15679 (W14282, W14289, W14288, W4844);
and G15680 (W14283, W15447, W4840);
and G15681 (W14284, W15447, W15446, W14286);
nand G15682 (W14285, W4804, W12618);
not G15683 (W14286, W4844);
not G15684 (W14287, W14289);
not G15685 (W14288, W4840);
not G15686 (W14289, W15055);
not G15687 (W14290, W4848);
nand G15688 (W14291, W4804, W12618);
and G15689 (W14292, W14287, W4844, W14290);
and G15690 (W14293, W14289, W4844, W4848);
and G15691 (W14294, W15448, W14289, W14290);
and G15692 (W14295, W15448, W14287, W4848);
nand G15693 (W14296, W4804, W12618);
nand G15694 (W14297, W14286, W14288);
nand G15695 (W14298, W4804, W12618);
nand G15696 (W14299, W4804, W12617);
nand G15697 (W14300, W4804, W12616);
nand G15698 (W14301, W4804, W12617);
nand G15699 (W14302, W4804, W12616);
nand G15700 (W14303, W4804, W12617);
nand G15701 (W14304, W4804, W12616);
nand G15702 (W14305, W4804, W12617);
nand G15703 (W14306, W4804, W12616);
nand G15704 (W14307, W15449, W15450);
nand G15705 (W14308, W15370, W15450);
nor G15706 (W14309, W15451, W15452, W15453);
nor G15707 (W14310, W15454, W15455, W15456);
and G15708 (W14311, W15454, W15455, W15456);
nand G15709 (W14312, W15457, W12616);
nand G15710 (W14313, W15457, W12617);
nand G15711 (W14314, W15457, W12618);
nand G15712 (W14315, W15458, W15459);
nand G15713 (W14316, W15460, W15461);
nand G15714 (W14317, W4835, W15461);
nand G15715 (W14318, W15462, W15463);
nand G15716 (W14319, W15464, W15463);
nor G15717 (W14320, W12594, W15465, W15466, W15467);
nand G15718 (W14321, W15468, W12616);
nand G15719 (W14322, W15468, W12617);
nand G15720 (W14323, W15468, W12618);
not G15721 (W14324, I95);
not G15722 (W14325, I94);
not G15723 (W14326, I1456);
nand G15724 (W14327, W15469, W9880);
nand G15725 (W14328, W15469, W9880);
nand G15726 (W14329, W15469, W9880);
nand G15727 (W14330, W15469, W9880);
nand G15728 (W14331, W15469, W9880);
nand G15729 (W14332, W15469, W9880);
and G15730 (W14333, W14244, W9918);
and G15731 (W14334, W14245, W9915);
and G15732 (W14335, W9880, W9912);
nand G15733 (W14336, W15469, W9880);
nand G15734 (W14337, W15469, W9880);
and G15735 (W14338, W14244, W9927);
and G15736 (W14339, W14245, W9924);
and G15737 (W14340, W9880, W9921);
nand G15738 (W14341, W15469, W9880);
nand G15739 (W14342, W15469, W9880);
nand G15740 (W14343, W15469, W14245);
nand G15741 (W14344, W15469, W14244);
nand G15742 (W14345, W15469, W14245);
nand G15743 (W14346, W15469, W14244);
nand G15744 (W14347, W15469, W14245);
nand G15745 (W14348, W15469, W14244);
nand G15746 (W14349, W15469, W14245);
nand G15747 (W14350, W15469, W14244);
nand G15748 (W14351, W15469, W14245);
nand G15749 (W14352, W15469, W14244);
nand G15750 (W14353, W15469, W14245);
nand G15751 (W14354, W15469, W14244);
nand G15752 (W14355, W15469, W14245);
nand G15753 (W14356, W15469, W14245);
nand G15754 (W14357, W15469, W14244);
nand G15755 (W14358, W15469, W14245);
nand G15756 (W14359, W15469, W14244);
nand G15757 (W14360, W15469, W14245);
nand G15758 (W14361, W15469, W14244);
nand G15759 (W14362, W15469, W14244);
not G15760 (W14363, W15470);
not G15761 (W14364, W15471);
not G15762 (W14365, W15472);
not G15763 (W14366, W15473);
not G15764 (W14367, W15474);
not G15765 (W14368, W15475);
not G15766 (W14369, W15476);
not G15767 (W14370, W15477);
not G15768 (W14371, W15478);
not G15769 (W14372, W15479);
nand G15770 (W14373, W15480, W9880);
nand G15771 (W14374, W15480, W14245);
nand G15772 (W14375, W15480, W14244);
nand G15773 (W14376, W15480, W9880);
nand G15774 (W14377, W15480, W14245);
nand G15775 (W14378, W15480, W14244);
nand G15776 (W14379, W15480, W9880);
nand G15777 (W14380, W15480, W14245);
nand G15778 (W14381, W15480, W14244);
nand G15779 (W14382, W15480, W9880);
nand G15780 (W14383, W15480, W14245);
nand G15781 (W14384, W15480, W14244);
nor G15782 (W14385, W15481, W15482);
not G15783 (W14386, W15483);
and G15784 (W14387, W15484, W15485);
and G15785 (W14388, W15486, W15487);
not G15786 (W14389, W14406);
and G15787 (W14390, W15488, W15489);
and G15788 (W14391, W15490, W15491);
not G15789 (W14392, W14406);
nor G15790 (W14393, W15481, W15492);
and G15791 (W14394, W15493, W15494);
and G15792 (W14395, W15495, W15496);
not G15793 (W14396, W14406);
and G15794 (W14397, W15497, W15498);
and G15795 (W14398, W15499, W15500);
not G15796 (W14399, W14406);
nor G15797 (W14400, W15501, W15481, W15502);
and G15798 (W14401, W15503, W15504);
and G15799 (W14402, W15505, W15506);
not G15800 (W14403, W14406);
nor G15801 (W14404, W15507, W15481);
not G15802 (W14405, W15508);
not G15803 (W14406, W15509);
nand G15804 (W14407, W14411, W15510);
nand G15805 (W14408, W14400, W15510);
nand G15806 (W14409, W15511, W15512);
nand G15807 (W14410, W15513, W15512);
nor G15808 (W14411, W15501, W15481, W15514);
and G15809 (W14412, W15515, W15516);
and G15810 (W14413, W15517, W15518);
not G15811 (W14414, W14406);
not G15812 (W14415, W15481);
and G15813 (W14416, W15519, W15520);
and G15814 (W14417, W15521, W15522);
not G15815 (W14418, W14406);
and G15816 (W14419, W15523, W15524);
and G15817 (W14420, W15525, W15526);
not G15818 (W14421, W14406);
nand G15819 (W14422, W15527, W13641);
nand G15820 (W14423, W15527, W10090);
nand G15821 (W14424, W15527, W15528);
not G15822 (W14425, W15529);
not G15823 (W14426, W15530);
and G15824 (W14427, W15531, W15532);
nand G15825 (W14428, W15533, W13641);
nand G15826 (W14429, W15533, W10090);
nand G15827 (W14430, W15533, W15528);
nand G15828 (W14431, W9958, W13641);
nand G15829 (W14432, W9958, W10090);
nand G15830 (W14433, W9958, W15528);
nand G15831 (W14434, W9958, W13641);
nand G15832 (W14435, W9958, W10090);
nand G15833 (W14436, W9958, W15528);
nand G15834 (W14437, W15533, W13641);
nand G15835 (W14438, W15533, W10090);
nand G15836 (W14439, W15533, W15528);
nand G15837 (W14440, W15533, W13641);
nand G15838 (W14441, W15533, W10090);
nand G15839 (W14442, W15533, W15528);
nand G15840 (W14443, W15533, W13641);
nand G15841 (W14444, W15533, W10090);
nand G15842 (W14445, W15533, W15528);
nand G15843 (W14446, W15533, W13641);
nand G15844 (W14447, W15533, W10090);
nand G15845 (W14448, W15533, W15528);
nand G15846 (W14449, W15533, W13641);
nand G15847 (W14450, W15533, W10090);
nand G15848 (W14451, W15533, W15528);
nand G15849 (W14452, W15533, W13641);
nand G15850 (W14453, W15533, W10090);
nand G15851 (W14454, W15533, W15528);
nand G15852 (W14455, W15533, W13641);
nand G15853 (W14456, W15533, W10090);
nand G15854 (W14457, W15533, W15528);
nand G15855 (W14458, W15533, W13641);
nand G15856 (W14459, W15533, W10090);
nand G15857 (W14460, W15533, W15528);
nand G15858 (W14461, W15533, W13641);
nand G15859 (W14462, W15533, W10090);
nand G15860 (W14463, W15533, W15528);
nand G15861 (W14464, W15533, W13641);
nand G15862 (W14465, W15533, W10090);
nand G15863 (W14466, W15533, W15528);
not G15864 (W14467, W15534);
not G15865 (W14468, W15535);
not G15866 (W14469, W15536);
not G15867 (W14470, W15537);
not G15868 (W14471, W15538);
not G15869 (W14472, W15539);
not G15870 (W14473, W15540);
not G15871 (W14474, W15541);
not G15872 (W14475, W15542);
not G15873 (W14476, W15543);
not G15874 (W14477, W14479);
not G15875 (W14478, W15544);
not G15876 (W14479, W15545);
not G15877 (W14480, W15546);
not G15878 (W14481, W14483);
not G15879 (W14482, W15547);
not G15880 (W14483, W15548);
not G15881 (W14484, W14486);
not G15882 (W14485, W15549);
not G15883 (W14486, W15550);
not G15884 (W14487, W14489);
not G15885 (W14488, W15551);
not G15886 (W14489, W15552);
not G15887 (W14490, W14492);
not G15888 (W14491, W15553);
not G15889 (W14492, W15554);
nand G15890 (W14493, W15555, W15556);
not G15891 (W14494, I1457);
not G15892 (W14495, I221);
not G15893 (W14496, W14497);
not G15894 (W14497, W15557);
not G15895 (W14498, W4985);
not G15896 (W14499, W15558);
not G15897 (W14500, W15559);
not G15898 (W14501, W15560);
not G15899 (W14502, W15561);
not G15900 (W14503, W15562);
not G15901 (W14504, W12973);
not G15902 (W14505, W15563);
not G15903 (W14506, W15564);
not G15904 (W14507, W14509);
not G15905 (W14508, W15565);
not G15906 (W14509, W15566);
not G15907 (W14510, I1458);
not G15908 (W14511, W15567);
not G15909 (W14512, W14514);
not G15910 (W14513, W15568);
not G15911 (W14514, W15569);
not G15912 (W14515, W14517);
not G15913 (W14516, W15570);
not G15914 (W14517, W15571);
not G15915 (W14518, W14520);
not G15916 (W14519, W15572);
not G15917 (W14520, W15573);
not G15918 (W14521, W14523);
not G15919 (W14522, W15574);
not G15920 (W14523, W15575);
not G15921 (W14524, W14526);
not G15922 (W14525, W15576);
not G15923 (W14526, W15577);
not G15924 (W14527, W14529);
not G15925 (W14528, I1459);
not G15926 (W14529, W15578);
not G15927 (W14530, W15579);
nand G15928 (W14531, W15580, W15581, W10654);
nand G15929 (W14532, W15582, W13022);
nand G15930 (W14533, W15582, W13023);
nand G15931 (W14534, W15582, W13024);
and G15932 (W14535, W15583, W15584);
and G15933 (W14536, W15585, W15586);
not G15934 (W14537, W15587);
not G15935 (W14538, W15588);
and G15936 (W14539, W15589, W15590);
and G15937 (W14540, W15591, W15592);
and G15938 (W14541, W15593, W15594);
and G15939 (W14542, W15595, W15596);
and G15940 (W14543, W15597, W15598);
and G15941 (W14544, W15599, W15600);
and G15942 (W14545, W15601, W15602);
and G15943 (W14546, W15603, W15604);
and G15944 (W14547, W15605, W15606);
and G15945 (W14548, W15607, W15608);
and G15946 (W14549, W15609, W15610);
and G15947 (W14550, W15611, W15612);
and G15948 (W14551, W15613, W15614);
and G15949 (W14552, W15615, W15616);
and G15950 (W14553, W15617, W15618);
and G15951 (W14554, W15619, W15620);
and G15952 (W14555, W15621, W15622);
and G15953 (W14556, W15623, W15624);
and G15954 (W14557, W14530, W12911);
nand G15955 (W14558, W15625, W15626);
not G15956 (W14559, W15627);
nand G15957 (W14560, W15628, W15629);
and G15958 (W14561, W14569, W15630);
and G15959 (W14562, W14570, W15631, W12911);
not G15960 (W14563, W15632);
nand G15961 (W14564, W15633, W13024);
nand G15962 (W14565, W15633, W13023);
nand G15963 (W14566, W15633, W13022);
or G15964 (W14567, W15634, W15635);
or G15965 (W14568, W10655, W15636);
not G15966 (W14569, W15637);
not G15967 (W14570, W15638);
not G15968 (W14571, W15632);
not G15969 (W14572, W15558);
and G15970 (W14573, W14580, W5111);
and G15971 (W14574, W14582, W15639, W5123);
and G15972 (W14575, W14582, W14581, W5119);
and G15973 (W14576, W15640, W5115);
and G15974 (W14577, W15640, W15639, W14579);
nand G15975 (W14578, W5079, W13024);
not G15976 (W14579, W5119);
not G15977 (W14580, W14582);
not G15978 (W14581, W5115);
not G15979 (W14582, W15055);
not G15980 (W14583, W5123);
nand G15981 (W14584, W5079, W13024);
and G15982 (W14585, W14580, W5119, W14583);
and G15983 (W14586, W14582, W5119, W5123);
and G15984 (W14587, W15641, W14582, W14583);
and G15985 (W14588, W15641, W14580, W5123);
nand G15986 (W14589, W5079, W13024);
nand G15987 (W14590, W14579, W14581);
nand G15988 (W14591, W5079, W13024);
nand G15989 (W14592, W5079, W13023);
nand G15990 (W14593, W5079, W13022);
nand G15991 (W14594, W5079, W13023);
nand G15992 (W14595, W5079, W13022);
nand G15993 (W14596, W5079, W13023);
nand G15994 (W14597, W5079, W13022);
nand G15995 (W14598, W5079, W13023);
nand G15996 (W14599, W5079, W13022);
nand G15997 (W14600, W15642, W15643);
nand G15998 (W14601, W15563, W15643);
nor G15999 (W14602, W15644, W15645, W15646);
nor G16000 (W14603, W15647, W15648, W15649);
and G16001 (W14604, W15647, W15648, W15649);
nand G16002 (W14605, W15650, W13022);
nand G16003 (W14606, W15650, W13023);
nand G16004 (W14607, W15650, W13024);
nand G16005 (W14608, W15651, W15652);
nand G16006 (W14609, W15653, W15654);
nand G16007 (W14610, W5110, W15654);
nand G16008 (W14611, W15655, W15656);
nand G16009 (W14612, W15657, W15656);
nor G16010 (W14613, W13000, W15658, W15659, W15660);
nand G16011 (W14614, W15661, W13022);
nand G16012 (W14615, W15661, W13023);
nand G16013 (W14616, W15661, W13024);
not G16014 (W14617, I144);
not G16015 (W14618, I143);
not G16016 (W14619, I1460);
nand G16017 (W14620, W15662, W10653);
nand G16018 (W14621, W15662, W10653);
nand G16019 (W14622, W15662, W10653);
nand G16020 (W14623, W15662, W10653);
nand G16021 (W14624, W15662, W10653);
and G16022 (W14625, W14537, W10691);
and G16023 (W14626, W14538, W10688);
and G16024 (W14627, W10653, W10685);
nand G16025 (W14628, W15662, W10653);
nand G16026 (W14629, W15662, W10653);
and G16027 (W14630, W14537, W10700);
and G16028 (W14631, W14538, W10697);
and G16029 (W14632, W10653, W10694);
nand G16030 (W14633, W15662, W10653);
nand G16031 (W14634, W15662, W10653);
nand G16032 (W14635, W15662, W14538);
nand G16033 (W14636, W15662, W14537);
nand G16034 (W14637, W15662, W14538);
nand G16035 (W14638, W15662, W14537);
nand G16036 (W14639, W15662, W14538);
nand G16037 (W14640, W15662, W14537);
nand G16038 (W14641, W15662, W14538);
nand G16039 (W14642, W15662, W14537);
nand G16040 (W14643, W15662, W14538);
nand G16041 (W14644, W15662, W14537);
nand G16042 (W14645, W15662, W14538);
nand G16043 (W14646, W15662, W14537);
nand G16044 (W14647, W15662, W14538);
nand G16045 (W14648, W15662, W14538);
nand G16046 (W14649, W15662, W14537);
nand G16047 (W14650, W15662, W14538);
nand G16048 (W14651, W15662, W14537);
nand G16049 (W14652, W15662, W14538);
nand G16050 (W14653, W15662, W14537);
nand G16051 (W14654, W15662, W14537);
nand G16052 (W14655, W15662, W10653);
not G16053 (W14656, W15663);
not G16054 (W14657, W15664);
not G16055 (W14658, W15665);
not G16056 (W14659, W15666);
not G16057 (W14660, W15667);
not G16058 (W14661, W15668);
not G16059 (W14662, W15669);
not G16060 (W14663, W15670);
not G16061 (W14664, W15671);
not G16062 (W14665, W15672);
nand G16063 (W14666, W15673, W10653);
nand G16064 (W14667, W15673, W14538);
nand G16065 (W14668, W15673, W14537);
nand G16066 (W14669, W15673, W10653);
nand G16067 (W14670, W15673, W14538);
nand G16068 (W14671, W15673, W14537);
nand G16069 (W14672, W15673, W10653);
nand G16070 (W14673, W15673, W14538);
nand G16071 (W14674, W15673, W14537);
nand G16072 (W14675, W15673, W10653);
nand G16073 (W14676, W15673, W14538);
nand G16074 (W14677, W15673, W14537);
nor G16075 (W14678, W15674, W15675);
not G16076 (W14679, W15676);
and G16077 (W14680, W15677, W15678);
and G16078 (W14681, W15679, W15680);
not G16079 (W14682, W14699);
and G16080 (W14683, W15681, W15682);
and G16081 (W14684, W15683, W15684);
not G16082 (W14685, W14699);
nor G16083 (W14686, W15674, W15685);
and G16084 (W14687, W15686, W15687);
and G16085 (W14688, W15688, W15689);
not G16086 (W14689, W14699);
and G16087 (W14690, W15690, W15691);
and G16088 (W14691, W15692, W15693);
not G16089 (W14692, W14699);
nor G16090 (W14693, W15694, W15674, W15695);
and G16091 (W14694, W15696, W15697);
and G16092 (W14695, W15698, W15699);
not G16093 (W14696, W14699);
nor G16094 (W14697, W15700, W15674);
not G16095 (W14698, W15701);
not G16096 (W14699, W15702);
nand G16097 (W14700, W14704, W15703);
nand G16098 (W14701, W14693, W15703);
nand G16099 (W14702, W15704, W15705);
nand G16100 (W14703, W15706, W15705);
nor G16101 (W14704, W15694, W15674, W15707);
and G16102 (W14705, W15708, W15709);
and G16103 (W14706, W15710, W15711);
not G16104 (W14707, W14699);
not G16105 (W14708, W15674);
and G16106 (W14709, W15712, W15713);
and G16107 (W14710, W15714, W15715);
not G16108 (W14711, W14699);
and G16109 (W14712, W15716, W15717);
and G16110 (W14713, W15718, W15719);
not G16111 (W14714, W14699);
nand G16112 (W14715, W15720, W13640);
nand G16113 (W14716, W15720, W10863);
nand G16114 (W14717, W15720, W15721);
not G16115 (W14718, W15722);
not G16116 (W14719, W15723);
and G16117 (W14720, W15724, W15725);
nand G16118 (W14721, W15726, W13640);
nand G16119 (W14722, W15726, W10863);
nand G16120 (W14723, W15726, W15721);
nand G16121 (W14724, W10731, W13640);
nand G16122 (W14725, W10731, W10863);
nand G16123 (W14726, W10731, W15721);
nand G16124 (W14727, W10731, W13640);
nand G16125 (W14728, W10731, W10863);
nand G16126 (W14729, W10731, W15721);
nand G16127 (W14730, W15726, W13640);
nand G16128 (W14731, W15726, W10863);
nand G16129 (W14732, W15726, W15721);
nand G16130 (W14733, W15726, W13640);
nand G16131 (W14734, W15726, W10863);
nand G16132 (W14735, W15726, W15721);
nand G16133 (W14736, W15726, W13640);
nand G16134 (W14737, W15726, W10863);
nand G16135 (W14738, W15726, W15721);
nand G16136 (W14739, W15726, W13640);
nand G16137 (W14740, W15726, W10863);
nand G16138 (W14741, W15726, W15721);
nand G16139 (W14742, W15726, W13640);
nand G16140 (W14743, W15726, W10863);
nand G16141 (W14744, W15726, W15721);
nand G16142 (W14745, W15726, W13640);
nand G16143 (W14746, W15726, W10863);
nand G16144 (W14747, W15726, W15721);
nand G16145 (W14748, W15726, W13640);
nand G16146 (W14749, W15726, W10863);
nand G16147 (W14750, W15726, W15721);
nand G16148 (W14751, W15726, W13640);
nand G16149 (W14752, W15726, W10863);
nand G16150 (W14753, W15726, W15721);
nand G16151 (W14754, W15726, W13640);
nand G16152 (W14755, W15726, W10863);
nand G16153 (W14756, W15726, W15721);
nand G16154 (W14757, W15726, W13640);
nand G16155 (W14758, W15726, W10863);
nand G16156 (W14759, W15726, W15721);
not G16157 (W14760, W15727);
not G16158 (W14761, W15728);
not G16159 (W14762, W15729);
not G16160 (W14763, W15730);
not G16161 (W14764, W15731);
not G16162 (W14765, W15732);
not G16163 (W14766, W15733);
not G16164 (W14767, W15734);
not G16165 (W14768, W15735);
not G16166 (W14769, W15736);
not G16167 (W14770, W15737);
not G16168 (W14771, W15737);
not G16169 (W14772, W15738);
not G16170 (W14773, W15739);
not G16171 (W14774, W15740);
not G16172 (W14775, W15741);
not G16173 (W14776, W15742);
nand G16174 (W14777, W15743, W15744);
not G16175 (W14778, I1461);
not G16176 (W14779, I222);
not G16177 (W14780, W15745);
not G16178 (W14781, W5260);
not G16179 (W14782, W15746);
not G16180 (W14783, W15747);
not G16181 (W14784, W15748);
not G16182 (W14785, W15749);
not G16183 (W14786, W15750);
not G16184 (W14787, W13368);
not G16185 (W14788, W15751);
not G16186 (W14789, W15752);
not G16187 (W14790, W15753);
not G16188 (W14791, I1462);
not G16189 (W14792, W15754);
not G16190 (W14793, W15755);
not G16191 (W14794, W15756);
not G16192 (W14795, W15757);
not G16193 (W14796, W15758);
not G16194 (W14797, W15759);
not G16195 (W14798, W14800);
not G16196 (W14799, I1463);
not G16197 (W14800, W15760);
not G16198 (W14801, W15761);
nand G16199 (W14802, W15762, W15763, W11427);
nand G16200 (W14803, W15764, W13417);
nand G16201 (W14804, W15764, W13418);
nand G16202 (W14805, W15764, W13419);
and G16203 (W14806, W15765, W15766);
and G16204 (W14807, W15767, W15768);
not G16205 (W14808, W15769);
not G16206 (W14809, W15770);
and G16207 (W14810, W15771, W15772);
and G16208 (W14811, W15773, W15774);
and G16209 (W14812, W15775, W15776);
and G16210 (W14813, W15777, W15778);
and G16211 (W14814, W15779, W15780);
and G16212 (W14815, W15781, W15782);
and G16213 (W14816, W15783, W15784);
and G16214 (W14817, W15785, W15786);
and G16215 (W14818, W15787, W15788);
and G16216 (W14819, W15789, W15790);
and G16217 (W14820, W15791, W15792);
and G16218 (W14821, W15793, W15794);
and G16219 (W14822, W15795, W15796);
and G16220 (W14823, W15797, W15798);
and G16221 (W14824, W15799, W15800);
and G16222 (W14825, W15801, W15802);
and G16223 (W14826, W15803, W15804);
and G16224 (W14827, W15805, W15806);
and G16225 (W14828, W14801, W13306);
nand G16226 (W14829, W15807, W15808);
not G16227 (W14830, W15809);
nand G16228 (W14831, W15810, W15811);
and G16229 (W14832, W14840, W15812);
and G16230 (W14833, W14841, W15813, W13306);
not G16231 (W14834, W15814);
nand G16232 (W14835, W15815, W13419);
nand G16233 (W14836, W15815, W13418);
nand G16234 (W14837, W15815, W13417);
or G16235 (W14838, W15816, W15817);
or G16236 (W14839, W11428, W15818);
not G16237 (W14840, W15819);
not G16238 (W14841, W15820);
not G16239 (W14842, W15814);
not G16240 (W14843, W15746);
and G16241 (W14844, W14851, W5386);
and G16242 (W14845, W14853, W15821, W5398);
and G16243 (W14846, W14853, W14852, W5394);
and G16244 (W14847, W15822, W5390);
and G16245 (W14848, W15822, W15821, W14850);
nand G16246 (W14849, W5354, W13419);
not G16247 (W14850, W5394);
not G16248 (W14851, W14853);
not G16249 (W14852, W5390);
not G16250 (W14853, W15055);
not G16251 (W14854, W5398);
nand G16252 (W14855, W5354, W13419);
and G16253 (W14856, W14851, W5394, W14854);
and G16254 (W14857, W14853, W5394, W5398);
and G16255 (W14858, W15823, W14853, W14854);
and G16256 (W14859, W15823, W14851, W5398);
nand G16257 (W14860, W5354, W13419);
nand G16258 (W14861, W14850, W14852);
nand G16259 (W14862, W5354, W13419);
nand G16260 (W14863, W5354, W13418);
nand G16261 (W14864, W5354, W13417);
nand G16262 (W14865, W5354, W13418);
nand G16263 (W14866, W5354, W13417);
nand G16264 (W14867, W5354, W13418);
nand G16265 (W14868, W5354, W13417);
nand G16266 (W14869, W5354, W13418);
nand G16267 (W14870, W5354, W13417);
nand G16268 (W14871, W15824, W15825);
nand G16269 (W14872, W15751, W15825);
nor G16270 (W14873, W15826, W15827, W15828);
nor G16271 (W14874, W15829, W15830, W15831);
and G16272 (W14875, W15829, W15830, W15831);
nand G16273 (W14876, W15832, W13417);
nand G16274 (W14877, W15832, W13418);
nand G16275 (W14878, W15832, W13419);
nand G16276 (W14879, W15833, W15834);
nand G16277 (W14880, W15835, W15836);
nand G16278 (W14881, W5385, W15836);
nand G16279 (W14882, W15837, W15838);
nand G16280 (W14883, W15839, W15838);
nor G16281 (W14884, W13395, W15840, W15841, W15842);
nand G16282 (W14885, W15843, W13417);
nand G16283 (W14886, W15843, W13418);
nand G16284 (W14887, W15843, W13419);
not G16285 (W14888, I193);
not G16286 (W14889, I192);
not G16287 (W14890, I1464);
nand G16288 (W14891, W15844, W11426);
nand G16289 (W14892, W15844, W11426);
nand G16290 (W14893, W15844, W11426);
nand G16291 (W14894, W15844, W11426);
and G16292 (W14895, W14808, W11464);
and G16293 (W14896, W14809, W11461);
and G16294 (W14897, W11426, W11458);
nand G16295 (W14898, W15844, W11426);
nand G16296 (W14899, W15844, W11426);
and G16297 (W14900, W14808, W11473);
and G16298 (W14901, W14809, W11470);
and G16299 (W14902, W11426, W11467);
nand G16300 (W14903, W15844, W11426);
nand G16301 (W14904, W15844, W11426);
nand G16302 (W14905, W15844, W14809);
nand G16303 (W14906, W15844, W14808);
nand G16304 (W14907, W15844, W14809);
nand G16305 (W14908, W15844, W14808);
nand G16306 (W14909, W15844, W14809);
nand G16307 (W14910, W15844, W14808);
nand G16308 (W14911, W15844, W14809);
nand G16309 (W14912, W15844, W14808);
nand G16310 (W14913, W15844, W14809);
nand G16311 (W14914, W15844, W14808);
nand G16312 (W14915, W15844, W14809);
nand G16313 (W14916, W15844, W14808);
nand G16314 (W14917, W15844, W14809);
nand G16315 (W14918, W15844, W14809);
nand G16316 (W14919, W15844, W14808);
nand G16317 (W14920, W15844, W14809);
nand G16318 (W14921, W15844, W14808);
nand G16319 (W14922, W15844, W14809);
nand G16320 (W14923, W15844, W14808);
nand G16321 (W14924, W15844, W14808);
nand G16322 (W14925, W15844, W11426);
nand G16323 (W14926, W15844, W11426);
not G16324 (W14927, W15845);
not G16325 (W14928, W15846);
not G16326 (W14929, W15847);
not G16327 (W14930, W15848);
not G16328 (W14931, W15849);
not G16329 (W14932, W15850);
not G16330 (W14933, W15851);
not G16331 (W14934, W15852);
not G16332 (W14935, W15853);
not G16333 (W14936, W15854);
nand G16334 (W14937, W15855, W11426);
nand G16335 (W14938, W15855, W14809);
nand G16336 (W14939, W15855, W14808);
nand G16337 (W14940, W15855, W11426);
nand G16338 (W14941, W15855, W14809);
nand G16339 (W14942, W15855, W14808);
nand G16340 (W14943, W15855, W11426);
nand G16341 (W14944, W15855, W14809);
nand G16342 (W14945, W15855, W14808);
nand G16343 (W14946, W15855, W11426);
nand G16344 (W14947, W15855, W14809);
nand G16345 (W14948, W15855, W14808);
not G16346 (W14949, W15856);
not G16347 (W14950, W15857);
nand G16348 (W14951, W11616, W14952);
nor G16349 (W14952, W11653, W15858);
not G16350 (W14953, W15859);
not G16351 (W14954, W15860);
nand G16352 (W14955, W11618, W14952);
not G16353 (W14956, W15861);
not G16354 (W14957, W15862);
not G16355 (W14958, W15863);
not G16356 (W14959, W15864);
nand G16357 (W14960, W15865, W15866);
nand G16358 (W14961, W14960, W14962);
nand G16359 (W14962, W15867, W15868);
nand G16360 (W14963, W15869, W15870);
nand G16361 (W14964, W14963, W14965);
nand G16362 (W14965, W15871, W15872);
and G16363 (W14966, W15873, I1391, W13575, W15874);
not G16364 (W14967, W15875);
not G16365 (W14968, W15876);
not G16366 (W14969, W15877);
not G16367 (W14970, W11644);
not G16368 (W14971, W15878);
not G16369 (W14972, W15879);
not G16370 (W14973, W15880);
not G16371 (W14974, W15881);
not G16372 (W14975, W15882);
not G16373 (W14976, W15883);
not G16374 (W14977, W14978);
not G16375 (W14978, W7899);
not G16376 (W14979, W15884);
not G16377 (W14980, W15885);
not G16378 (W14981, W15886);
nand G16379 (W14982, W15887, W15888);
nand G16380 (W14983, W15889, W15888);
nand G16381 (W14984, W15890, W15891);
nand G16382 (W14985, W15892, W15891);
not G16383 (W14986, W15893);
nand G16384 (W14987, W15894, W15895);
nand G16385 (W14988, W15896, W15895);
nand G16386 (W14989, W15897, W15898);
nand G16387 (W14990, W15899, W15898);
not G16388 (W14991, I451);
not G16389 (W14992, W15900);
not G16390 (W14993, W8244);
not G16391 (W14994, W14996);
nor G16392 (W14995, W15901, W15902);
not G16393 (W14996, W15903);
not G16394 (W14997, W11787);
not G16395 (W14998, W15000);
nor G16396 (W14999, W15904, W15905);
not G16397 (W15000, W15906);
not G16398 (W15001, W13607);
nor G16399 (W15002, W15907, W15908, W5289);
not G16400 (W15003, W15909);
nor G16401 (W15004, W15910, W5288, W15907);
not G16402 (W15005, W15911);
not G16403 (W15006, W8287);
not G16404 (W15007, W15009);
nor G16405 (W15008, W15912, W15913);
not G16406 (W15009, W15914);
not G16407 (W15010, W11814);
not G16408 (W15011, W15013);
nor G16409 (W15012, W15915, W15916);
not G16410 (W15013, W15917);
not G16411 (W15014, W13607);
nor G16412 (W15015, W15907, W15918, W5014);
not G16413 (W15016, W15919);
nor G16414 (W15017, W15920, W5013, W15907);
not G16415 (W15018, W15921);
not G16416 (W15019, W8330);
not G16417 (W15020, W15022);
nor G16418 (W15021, W15922, W15923);
not G16419 (W15022, W15924);
not G16420 (W15023, W11840);
not G16421 (W15024, W15026);
nor G16422 (W15025, W15925, W15926);
not G16423 (W15026, W15927);
not G16424 (W15027, W13607);
nor G16425 (W15028, W15907, W15928, W4739);
not G16426 (W15029, W15929);
nor G16427 (W15030, W15930, W4738, W15907);
not G16428 (W15031, W15931);
not G16429 (W15032, W8373);
not G16430 (W15033, W15035);
nor G16431 (W15034, W15932, W15933);
not G16432 (W15035, W15934);
not G16433 (W15036, W11866);
not G16434 (W15037, W15039);
nor G16435 (W15038, W15935, W15936);
not G16436 (W15039, W15937);
not G16437 (W15040, W13607);
nor G16438 (W15041, W15907, W15938, W4464);
not G16439 (W15042, W15939);
nor G16440 (W15043, W15940, W4463, W15907);
not G16441 (W15044, W15941);
nand G16442 (W15045, W15047, I502);
nand G16443 (W15046, W11874, I503);
nor G16444 (W15047, W15046, W11752);
not G16445 (W15048, I1465);
not G16446 (W15049, I1466);
not G16447 (W15050, I1467);
not G16448 (W15051, I1468);
not G16449 (W15052, W5250);
nor G16450 (W15053, W13654, W13653);
not G16451 (W15054, W15942);
not G16452 (W15055, W15943);
nor G16453 (W15056, W5252, W5250);
and G16454 (W15057, W11015, I455);
and G16455 (W15058, W11016, I456);
and G16456 (W15059, W11017, I457);
and G16457 (W15060, W11882, W11884, W11888);
not G16458 (W15061, W4975);
nor G16459 (W15062, W13689, W13688);
not G16460 (W15063, W15944);
nor G16461 (W15064, W4977, W4975);
and G16462 (W15065, W10242, I467);
and G16463 (W15066, W10243, I468);
and G16464 (W15067, W10244, I469);
not G16465 (W15068, W4700);
nor G16466 (W15069, W13723, W13722);
not G16467 (W15070, W15945);
nor G16468 (W15071, W4702, W4700);
and G16469 (W15072, W9469, I479);
and G16470 (W15073, W9470, I480);
and G16471 (W15074, W9471, I481);
not G16472 (W15075, W4425);
nor G16473 (W15076, W13757, W13756);
not G16474 (W15077, W15946);
nor G16475 (W15078, W4427, W4425);
and G16476 (W15079, W8696, I491);
and G16477 (W15080, W8697, I492);
and G16478 (W15081, W8698, I493);
nor G16479 (W15082, W15089, W11890);
and G16480 (W15083, W13785, I1396, W11882, I558);
not G16481 (W15084, W13783);
not G16482 (W15085, W15947);
nor G16483 (W15086, W15947, W13787);
nand G16484 (W15087, W15086, I557);
nor G16485 (W15088, W15087, W11884);
nand G16486 (W15089, W15088, I559);
not G16487 (W15090, W15948);
not G16488 (W15091, W15949);
not G16489 (W15092, W15102);
nor G16490 (W15093, W15950, W15951);
nor G16491 (W15094, W15111, W15091, W15952);
not G16492 (W15095, W15097);
nor G16493 (W15096, W15091, I1469);
not G16494 (W15097, W15953);
nor G16495 (W15098, W15111, W15091, W15954);
not G16496 (W15099, W15101);
nor G16497 (W15100, W15091, I1470);
not G16498 (W15101, W15955);
nand G16499 (W15102, I219, W15956);
nor G16500 (W15103, W15111, W15091, W15957);
not G16501 (W15104, W15106);
nor G16502 (W15105, W15091, I1471);
not G16503 (W15106, W15958);
nor G16504 (W15107, W15111, W15091, W15959);
not G16505 (W15108, W15110);
nor G16506 (W15109, W15091, I1472);
not G16507 (W15110, W15960);
not G16508 (W15111, I219);
not G16509 (W15112, W15961);
nor G16510 (W15113, W15111, W15091, W15962);
not G16511 (W15114, W15116);
nor G16512 (W15115, W15091, I1473);
not G16513 (W15116, W15963);
or G16514 (W15117, W15964, W15965);
not G16515 (W15118, W15966);
not G16516 (W15119, W15951);
nand G16517 (W15120, W13821, W13810);
nand G16518 (W15121, W15967, W15968);
nand G16519 (W15122, W15121, W15123);
nand G16520 (W15123, W15969, W15970);
not G16521 (W15124, W15971);
nor G16522 (W15125, W15111, W15091, W15972);
not G16523 (W15126, W15128);
nor G16524 (W15127, W15091, I1474);
not G16525 (W15128, W15973);
nor G16526 (W15129, W15111, W15091, W15974);
not G16527 (W15130, W15132);
nor G16528 (W15131, W15091, I1475);
not G16529 (W15132, W15975);
nor G16530 (W15133, W15111, W15091, W15976);
not G16531 (W15134, W15136);
nor G16532 (W15135, W15091, I1476);
not G16533 (W15136, W15977);
or G16534 (W15137, W15143, W8412);
not G16535 (W15138, W15978);
nor G16536 (W15139, W15979, W15980, W15981);
nor G16537 (W15140, W15982, W15983, W15984);
and G16538 (W15141, W15985, W15986, W15987);
and G16539 (W15142, W15988, W15989, W15990);
and G16540 (W15143, W8197, W15991, I1477);
nor G16541 (W15144, W15145, W11982);
nand G16542 (W15145, W15146, I262);
nor G16543 (W15146, W15147, W11988);
nand G16544 (W15147, W15148, I264);
nor G16545 (W15148, W15149, W11994);
nand G16546 (W15149, W15150, I266);
nor G16547 (W15150, W15151, W12000);
nand G16548 (W15151, W15152, I268);
nor G16549 (W15152, W15153, W12006);
nand G16550 (W15153, W8197, W13643);
not G16551 (W15154, W4692);
not G16552 (W15155, W8697);
not G16553 (W15156, I1478);
not G16554 (W15157, W4693);
not G16555 (W15158, W8697);
not G16556 (W15159, W4694);
not G16557 (W15160, W8697);
not G16558 (W15161, W4695);
not G16559 (W15162, W8697);
not G16560 (W15163, W4696);
not G16561 (W15164, W8697);
nand G16562 (W15165, W15992, W15993);
nand G16563 (W15166, W8372, W15993);
not G16564 (W15167, I199);
not G16565 (W15168, I198);
not G16566 (W15169, I1479);
not G16567 (W15170, W8696);
nor G16568 (W15171, W15244, W15994, W13984);
not G16569 (W15172, I1480);
not G16570 (W15173, I10);
not G16571 (W15174, I11);
nor G16572 (W15175, W13982, W15994, W12156);
not G16573 (W15176, W15995);
not G16574 (W15177, I1451);
not G16575 (W15178, W4742);
not G16576 (W15179, W12211);
not G16577 (W15180, I1481);
not G16578 (W15181, W4743);
not G16579 (W15182, W12211);
not G16580 (W15183, W4744);
not G16581 (W15184, W12211);
not G16582 (W15185, W4745);
not G16583 (W15186, W12211);
not G16584 (W15187, W4746);
not G16585 (W15188, W12211);
not G16586 (W15189, W4747);
not G16587 (W15190, W12211);
not G16588 (W15191, W13996);
nor G16589 (W15192, W15996, W15997, W15998);
nor G16590 (W15193, W15999, W16000);
not G16591 (W15194, W16001);
not G16592 (W15195, W16002);
nor G16593 (W15196, W16003, W16004);
not G16594 (W15197, W15199);
nand G16595 (W15198, W9021, W16005);
not G16596 (W15199, W16006);
not G16597 (W15200, I50);
not G16598 (W15201, I49);
nor G16599 (W15202, W16007, W16008);
not G16600 (W15203, W15205);
nor G16601 (W15204, W16009, W16010);
not G16602 (W15205, W16011);
nor G16603 (W15206, W16012, W16013);
not G16604 (W15207, W15209);
nor G16605 (W15208, W16014, W16015);
not G16606 (W15209, W16016);
nor G16607 (W15210, W16017, W16018);
not G16608 (W15211, W15213);
nor G16609 (W15212, W16019, W16020);
not G16610 (W15213, W16021);
nor G16611 (W15214, W16022, W16023);
not G16612 (W15215, W15217);
nand G16613 (W15216, W9017, W16005);
not G16614 (W15217, W16024);
nor G16615 (W15218, W16025, W16026);
not G16616 (W15219, W15221);
nand G16617 (W15220, W9025, W16005);
not G16618 (W15221, W16027);
nor G16619 (W15222, W16028, W16029);
not G16620 (W15223, W15225);
nand G16621 (W15224, W9033, W16005);
not G16622 (W15225, W16030);
nor G16623 (W15226, W16031, W16032);
not G16624 (W15227, W15229);
nor G16625 (W15228, W16033, W16034);
not G16626 (W15229, W16035);
nor G16627 (W15230, W16036, W16037);
not G16628 (W15231, W15233);
nor G16629 (W15232, W16038, W16039);
not G16630 (W15233, W16040);
nor G16631 (W15234, W16041, W16042);
not G16632 (W15235, W15237);
nand G16633 (W15236, W9013, W16005);
not G16634 (W15237, W16043);
nand G16635 (W15238, W16044, W16045);
nand G16636 (W15239, W13984, W16045);
nand G16637 (W15240, W16046, W16047);
nand G16638 (W15241, W16048, W16049);
nand G16639 (W15242, W15994, W16049);
not G16640 (W15243, W16050);
not G16641 (W15244, W16051);
nor G16642 (W15245, W16052, W16053, W16054);
nor G16643 (W15246, W16055, W16056);
not G16644 (W15247, W16057);
not G16645 (W15248, W16058);
nand G16646 (W15249, W16059, W16060, W16061);
not G16647 (W15250, W16051);
not G16648 (W15251, W16062);
not G16649 (W15252, W15874);
not G16650 (W15253, W4561);
nor G16651 (W15254, W13997, W13996);
nor G16652 (W15255, W4569, W4561);
nor G16653 (W15256, W12190, W16063, W12188);
nand G16654 (W15257, W15256, W15176);
and G16655 (W15258, W12210, W8942);
and G16656 (W15259, W12211, W8945);
and G16657 (W15260, W12212, W8948);
not G16658 (W15261, W16064);
not G16659 (W15262, W15176);
not G16660 (W15263, W16065);
or G16661 (W15264, W16066, W8940);
nand G16662 (W15265, W16067, W16068);
nand G16663 (W15266, W15263, W16068);
nor G16664 (W15267, W12188, W16069);
nand G16665 (W15268, W15267, W4560);
nor G16666 (W15269, W12188, W16070);
nand G16667 (W15270, W15269, W15271);
not G16668 (W15271, W16071);
nor G16669 (W15272, W16072, W16073);
not G16670 (W15273, W15271);
not G16671 (W15274, W16074);
or G16672 (W15275, W16075, W14027);
not G16673 (W15276, W16076);
nor G16674 (W15277, W16077, W9109);
nand G16675 (W15278, W15277, I740);
nor G16676 (W15279, W15278, W12259);
nand G16677 (W15280, W15279, I742);
nor G16678 (W15281, W15280, W12265);
nand G16679 (W15282, W15281, I744);
nor G16680 (W15283, W15282, W12271);
nand G16681 (W15284, W15283, I746);
nor G16682 (W15285, W15284, W12277);
nand G16683 (W15286, W15285, I748);
not G16684 (W15287, W16078);
not G16685 (W15288, W16079);
not G16686 (W15289, W15299);
nor G16687 (W15290, W16080, W16081);
nor G16688 (W15291, W15308, W15288, W16082);
not G16689 (W15292, W15294);
nor G16690 (W15293, W15288, I1482);
not G16691 (W15294, W16083);
nor G16692 (W15295, W15308, W15288, W16084);
not G16693 (W15296, W15298);
nor G16694 (W15297, W15288, I1483);
not G16695 (W15298, W16085);
nand G16696 (W15299, I220, W16086);
nor G16697 (W15300, W15308, W15288, W16087);
not G16698 (W15301, W15303);
nor G16699 (W15302, W15288, I1484);
not G16700 (W15303, W16088);
nor G16701 (W15304, W15308, W15288, W16089);
not G16702 (W15305, W15307);
nor G16703 (W15306, W15288, I1485);
not G16704 (W15307, W16090);
not G16705 (W15308, I220);
not G16706 (W15309, W16091);
nor G16707 (W15310, W15308, W15288, W16092);
not G16708 (W15311, W15313);
nor G16709 (W15312, W15288, I1486);
not G16710 (W15313, W16093);
or G16711 (W15314, W16094, W16095);
not G16712 (W15315, W16096);
not G16713 (W15316, W16081);
nand G16714 (W15317, W14118, W14107);
nand G16715 (W15318, W16097, W16098);
nand G16716 (W15319, W15318, W15320);
nand G16717 (W15320, W16099, W16100);
not G16718 (W15321, W16101);
nor G16719 (W15322, W15308, W15288, W16102);
not G16720 (W15323, W15325);
nor G16721 (W15324, W15288, I1487);
not G16722 (W15325, W16103);
nor G16723 (W15326, W15308, W15288, W16104);
not G16724 (W15327, W15329);
nor G16725 (W15328, W15288, I1488);
not G16726 (W15329, W16105);
nor G16727 (W15330, W15308, W15288, W16106);
not G16728 (W15331, W15333);
nor G16729 (W15332, W15288, I1489);
not G16730 (W15333, W16107);
or G16731 (W15334, W15340, W9185);
not G16732 (W15335, W16108);
nor G16733 (W15336, W16109, W16110, W16111);
nor G16734 (W15337, W16112, W16113, W16114);
and G16735 (W15338, W16115, W16116, W16117);
and G16736 (W15339, W16118, W16119, W16120);
and G16737 (W15340, W8193, W16121, I1490);
nor G16738 (W15341, W15342, W12388);
nand G16739 (W15342, W15343, I298);
nor G16740 (W15343, W15344, W12394);
nand G16741 (W15344, W15345, I300);
nor G16742 (W15345, W15346, W12400);
nand G16743 (W15346, W15347, I302);
nor G16744 (W15347, W15348, W12406);
nand G16745 (W15348, W15349, I304);
nor G16746 (W15349, W15350, W12412);
nand G16747 (W15350, W8193, W13642);
not G16748 (W15351, W4967);
not G16749 (W15352, W9470);
not G16750 (W15353, I1491);
not G16751 (W15354, W4968);
not G16752 (W15355, W9470);
not G16753 (W15356, W4969);
not G16754 (W15357, W9470);
not G16755 (W15358, W4970);
not G16756 (W15359, W9470);
not G16757 (W15360, W4971);
not G16758 (W15361, W9470);
nand G16759 (W15362, W16122, W16123);
nand G16760 (W15363, W8329, W16123);
not G16761 (W15364, W9469);
nor G16762 (W15365, W15438, W16124, W14278);
not G16763 (W15366, I1492);
not G16764 (W15367, I59);
not G16765 (W15368, I60);
nor G16766 (W15369, W14276, W16124, W12562);
not G16767 (W15370, W16125);
not G16768 (W15371, I1455);
not G16769 (W15372, W5017);
not G16770 (W15373, W12617);
not G16771 (W15374, I1493);
not G16772 (W15375, W5018);
not G16773 (W15376, W12617);
not G16774 (W15377, W5019);
not G16775 (W15378, W12617);
not G16776 (W15379, W5020);
not G16777 (W15380, W12617);
not G16778 (W15381, W5021);
not G16779 (W15382, W12617);
not G16780 (W15383, W5022);
not G16781 (W15384, W12617);
not G16782 (W15385, W14289);
nor G16783 (W15386, W16126, W16127, W16128);
nor G16784 (W15387, W16129, W16130);
not G16785 (W15388, W16131);
not G16786 (W15389, W16132);
nor G16787 (W15390, W16133, W16134);
not G16788 (W15391, W15393);
nand G16789 (W15392, W9794, W16135);
not G16790 (W15393, W16136);
not G16791 (W15394, I99);
not G16792 (W15395, I98);
nor G16793 (W15396, W16137, W16138);
not G16794 (W15397, W15399);
nor G16795 (W15398, W16139, W16140);
not G16796 (W15399, W16141);
nor G16797 (W15400, W16142, W16143);
not G16798 (W15401, W15403);
nor G16799 (W15402, W16144, W16145);
not G16800 (W15403, W16146);
nor G16801 (W15404, W16147, W16148);
not G16802 (W15405, W15407);
nor G16803 (W15406, W16149, W16150);
not G16804 (W15407, W16151);
nor G16805 (W15408, W16152, W16153);
not G16806 (W15409, W15411);
nand G16807 (W15410, W9790, W16135);
not G16808 (W15411, W16154);
nor G16809 (W15412, W16155, W16156);
not G16810 (W15413, W15415);
nand G16811 (W15414, W9798, W16135);
not G16812 (W15415, W16157);
nor G16813 (W15416, W16158, W16159);
not G16814 (W15417, W15419);
nand G16815 (W15418, W9806, W16135);
not G16816 (W15419, W16160);
nor G16817 (W15420, W16161, W16162);
not G16818 (W15421, W15423);
nor G16819 (W15422, W16163, W16164);
not G16820 (W15423, W16165);
nor G16821 (W15424, W16166, W16167);
not G16822 (W15425, W15427);
nor G16823 (W15426, W16168, W16169);
not G16824 (W15427, W16170);
nor G16825 (W15428, W16171, W16172);
not G16826 (W15429, W15431);
nand G16827 (W15430, W9786, W16135);
not G16828 (W15431, W16173);
nand G16829 (W15432, W16174, W16175);
nand G16830 (W15433, W14278, W16175);
nand G16831 (W15434, W16176, W16177);
nand G16832 (W15435, W16178, W16179);
nand G16833 (W15436, W16124, W16179);
not G16834 (W15437, W16180);
not G16835 (W15438, W16181);
nor G16836 (W15439, W16182, W16183, W16184);
nor G16837 (W15440, W16185, W16186);
not G16838 (W15441, W16187);
not G16839 (W15442, W16188);
nand G16840 (W15443, W16189, W16190, W16191);
not G16841 (W15444, W16181);
not G16842 (W15445, W16192);
not G16843 (W15446, W4836);
nor G16844 (W15447, W14290, W14289);
nor G16845 (W15448, W4844, W4836);
nor G16846 (W15449, W12596, W16193, W12594);
nand G16847 (W15450, W15449, W15370);
and G16848 (W15451, W12616, W9715);
and G16849 (W15452, W12617, W9718);
and G16850 (W15453, W12618, W9721);
not G16851 (W15454, W16194);
not G16852 (W15455, W15370);
not G16853 (W15456, W16195);
or G16854 (W15457, W16196, W9713);
nand G16855 (W15458, W16197, W16198);
nand G16856 (W15459, W15456, W16198);
nor G16857 (W15460, W12594, W16199);
nand G16858 (W15461, W15460, W4835);
nor G16859 (W15462, W12594, W16200);
nand G16860 (W15463, W15462, W15464);
not G16861 (W15464, W16201);
nor G16862 (W15465, W16202, W16203);
not G16863 (W15466, W15464);
not G16864 (W15467, W16204);
or G16865 (W15468, W16205, W14320);
not G16866 (W15469, W16206);
nor G16867 (W15470, W16207, W9882);
nand G16868 (W15471, W15470, I941);
nor G16869 (W15472, W15471, W12665);
nand G16870 (W15473, W15472, I943);
nor G16871 (W15474, W15473, W12671);
nand G16872 (W15475, W15474, I945);
nor G16873 (W15476, W15475, W12677);
nand G16874 (W15477, W15476, I947);
nor G16875 (W15478, W15477, W12683);
nand G16876 (W15479, W15478, I949);
not G16877 (W15480, W16208);
not G16878 (W15481, W16209);
not G16879 (W15482, W15492);
nor G16880 (W15483, W16210, W16211);
nor G16881 (W15484, W15501, W15481, W16212);
not G16882 (W15485, W15487);
nor G16883 (W15486, W15481, I1494);
not G16884 (W15487, W16213);
nor G16885 (W15488, W15501, W15481, W16214);
not G16886 (W15489, W15491);
nor G16887 (W15490, W15481, I1495);
not G16888 (W15491, W16215);
nand G16889 (W15492, I221, W16216);
nor G16890 (W15493, W15501, W15481, W16217);
not G16891 (W15494, W15496);
nor G16892 (W15495, W15481, I1496);
not G16893 (W15496, W16218);
nor G16894 (W15497, W15501, W15481, W16219);
not G16895 (W15498, W15500);
nor G16896 (W15499, W15481, I1497);
not G16897 (W15500, W16220);
not G16898 (W15501, I221);
not G16899 (W15502, W16221);
nor G16900 (W15503, W15501, W15481, W16222);
not G16901 (W15504, W15506);
nor G16902 (W15505, W15481, I1498);
not G16903 (W15506, W16223);
or G16904 (W15507, W16224, W16225);
not G16905 (W15508, W16226);
not G16906 (W15509, W16211);
nand G16907 (W15510, W14411, W14400);
nand G16908 (W15511, W16227, W16228);
nand G16909 (W15512, W15511, W15513);
nand G16910 (W15513, W16229, W16230);
not G16911 (W15514, W16231);
nor G16912 (W15515, W15501, W15481, W16232);
not G16913 (W15516, W15518);
nor G16914 (W15517, W15481, I1499);
not G16915 (W15518, W16233);
nor G16916 (W15519, W15501, W15481, W16234);
not G16917 (W15520, W15522);
nor G16918 (W15521, W15481, I1500);
not G16919 (W15522, W16235);
nor G16920 (W15523, W15501, W15481, W16236);
not G16921 (W15524, W15526);
nor G16922 (W15525, W15481, I1501);
not G16923 (W15526, W16237);
or G16924 (W15527, W15533, W9958);
not G16925 (W15528, W16238);
nor G16926 (W15529, W16239, W16240, W16241);
nor G16927 (W15530, W16242, W16243, W16244);
and G16928 (W15531, W16245, W16246, W16247);
and G16929 (W15532, W16248, W16249, W16250);
and G16930 (W15533, W8189, W16251, I1502);
nor G16931 (W15534, W15535, W12794);
nand G16932 (W15535, W15536, I334);
nor G16933 (W15536, W15537, W12800);
nand G16934 (W15537, W15538, I336);
nor G16935 (W15538, W15539, W12806);
nand G16936 (W15539, W15540, I338);
nor G16937 (W15540, W15541, W12812);
nand G16938 (W15541, W15542, I340);
nor G16939 (W15542, W15543, W12818);
nand G16940 (W15543, W8189, W13641);
not G16941 (W15544, W5242);
not G16942 (W15545, W10243);
not G16943 (W15546, I1503);
not G16944 (W15547, W5243);
not G16945 (W15548, W10243);
not G16946 (W15549, W5244);
not G16947 (W15550, W10243);
not G16948 (W15551, W5245);
not G16949 (W15552, W10243);
not G16950 (W15553, W5246);
not G16951 (W15554, W10243);
nand G16952 (W15555, W16252, W16253);
nand G16953 (W15556, W8286, W16253);
not G16954 (W15557, W10242);
nor G16955 (W15558, W15631, W16254, W14571);
not G16956 (W15559, I1504);
not G16957 (W15560, I108);
not G16958 (W15561, I109);
nor G16959 (W15562, W14569, W16254, W12968);
not G16960 (W15563, W16255);
not G16961 (W15564, I1459);
not G16962 (W15565, W5292);
not G16963 (W15566, W13023);
not G16964 (W15567, I1505);
not G16965 (W15568, W5293);
not G16966 (W15569, W13023);
not G16967 (W15570, W5294);
not G16968 (W15571, W13023);
not G16969 (W15572, W5295);
not G16970 (W15573, W13023);
not G16971 (W15574, W5296);
not G16972 (W15575, W13023);
not G16973 (W15576, W5297);
not G16974 (W15577, W13023);
not G16975 (W15578, W14582);
nor G16976 (W15579, W16256, W16257, W16258);
nor G16977 (W15580, W16259, W16260);
not G16978 (W15581, W16261);
not G16979 (W15582, W16262);
nor G16980 (W15583, W16263, W16264);
not G16981 (W15584, W15586);
nand G16982 (W15585, W10563, W16265);
not G16983 (W15586, W16266);
not G16984 (W15587, I148);
not G16985 (W15588, I147);
nor G16986 (W15589, W16267, W16268);
not G16987 (W15590, W15592);
nor G16988 (W15591, W16269, W16270);
not G16989 (W15592, W16271);
nor G16990 (W15593, W16272, W16273);
not G16991 (W15594, W15596);
nor G16992 (W15595, W16274, W16275);
not G16993 (W15596, W16276);
nor G16994 (W15597, W16277, W16278);
not G16995 (W15598, W15600);
nor G16996 (W15599, W16279, W16280);
not G16997 (W15600, W16281);
nor G16998 (W15601, W16282, W16283);
not G16999 (W15602, W15604);
nand G17000 (W15603, W10559, W16265);
not G17001 (W15604, W16284);
nor G17002 (W15605, W16285, W16286);
not G17003 (W15606, W15608);
nand G17004 (W15607, W10567, W16265);
not G17005 (W15608, W16287);
nor G17006 (W15609, W16288, W16289);
not G17007 (W15610, W15612);
nand G17008 (W15611, W10575, W16265);
not G17009 (W15612, W16290);
nor G17010 (W15613, W16291, W16292);
not G17011 (W15614, W15616);
nor G17012 (W15615, W16293, W16294);
not G17013 (W15616, W16295);
nor G17014 (W15617, W16296, W16297);
not G17015 (W15618, W15620);
nor G17016 (W15619, W16298, W16299);
not G17017 (W15620, W16300);
nor G17018 (W15621, W16301, W16302);
not G17019 (W15622, W15624);
nand G17020 (W15623, W10555, W16265);
not G17021 (W15624, W16303);
nand G17022 (W15625, W16304, W16305);
nand G17023 (W15626, W14571, W16305);
nand G17024 (W15627, W16306, W16307);
nand G17025 (W15628, W16308, W16309);
nand G17026 (W15629, W16254, W16309);
not G17027 (W15630, W16310);
not G17028 (W15631, W16311);
nor G17029 (W15632, W16312, W16313, W16314);
nor G17030 (W15633, W16315, W16316);
not G17031 (W15634, W16317);
not G17032 (W15635, W16318);
nand G17033 (W15636, W16319, W16320, W16321);
not G17034 (W15637, W16311);
not G17035 (W15638, W16322);
not G17036 (W15639, W5111);
nor G17037 (W15640, W14583, W14582);
nor G17038 (W15641, W5119, W5111);
nor G17039 (W15642, W13002, W16323, W13000);
nand G17040 (W15643, W15642, W15563);
and G17041 (W15644, W13022, W10488);
and G17042 (W15645, W13023, W10491);
and G17043 (W15646, W13024, W10494);
not G17044 (W15647, W16324);
not G17045 (W15648, W15563);
not G17046 (W15649, W16325);
or G17047 (W15650, W16326, W10486);
nand G17048 (W15651, W16327, W16328);
nand G17049 (W15652, W15649, W16328);
nor G17050 (W15653, W13000, W16329);
nand G17051 (W15654, W15653, W5110);
nor G17052 (W15655, W13000, W16330);
nand G17053 (W15656, W15655, W15657);
not G17054 (W15657, W16331);
nor G17055 (W15658, W16332, W16333);
not G17056 (W15659, W15657);
not G17057 (W15660, W16334);
or G17058 (W15661, W16335, W14613);
not G17059 (W15662, W16336);
nor G17060 (W15663, W16337, W10655);
nand G17061 (W15664, W15663, I1142);
nor G17062 (W15665, W15664, W13071);
nand G17063 (W15666, W15665, I1144);
nor G17064 (W15667, W15666, W13077);
nand G17065 (W15668, W15667, I1146);
nor G17066 (W15669, W15668, W13083);
nand G17067 (W15670, W15669, I1148);
nor G17068 (W15671, W15670, W13089);
nand G17069 (W15672, W15671, I1150);
not G17070 (W15673, W16338);
not G17071 (W15674, W16339);
not G17072 (W15675, W15685);
nor G17073 (W15676, W16340, W16341);
nor G17074 (W15677, W15694, W15674, W16342);
not G17075 (W15678, W15680);
nor G17076 (W15679, W15674, I1506);
not G17077 (W15680, W16343);
nor G17078 (W15681, W15694, W15674, W16344);
not G17079 (W15682, W15684);
nor G17080 (W15683, W15674, I1507);
not G17081 (W15684, W16345);
nand G17082 (W15685, I222, W16346);
nor G17083 (W15686, W15694, W15674, W16347);
not G17084 (W15687, W15689);
nor G17085 (W15688, W15674, I1508);
not G17086 (W15689, W16348);
nor G17087 (W15690, W15694, W15674, W16349);
not G17088 (W15691, W15693);
nor G17089 (W15692, W15674, I1509);
not G17090 (W15693, W16350);
not G17091 (W15694, I222);
not G17092 (W15695, W16351);
nor G17093 (W15696, W15694, W15674, W16352);
not G17094 (W15697, W15699);
nor G17095 (W15698, W15674, I1510);
not G17096 (W15699, W16353);
or G17097 (W15700, W16354, W16355);
not G17098 (W15701, W16356);
not G17099 (W15702, W16341);
nand G17100 (W15703, W14704, W14693);
nand G17101 (W15704, W16357, W16358);
nand G17102 (W15705, W15704, W15706);
nand G17103 (W15706, W16359, W16360);
not G17104 (W15707, W16361);
nor G17105 (W15708, W15694, W15674, W16362);
not G17106 (W15709, W15711);
nor G17107 (W15710, W15674, I1511);
not G17108 (W15711, W16363);
nor G17109 (W15712, W15694, W15674, W16364);
not G17110 (W15713, W15715);
nor G17111 (W15714, W15674, I1512);
not G17112 (W15715, W16365);
nor G17113 (W15716, W15694, W15674, W16366);
not G17114 (W15717, W15719);
nor G17115 (W15718, W15674, I1513);
not G17116 (W15719, W16367);
or G17117 (W15720, W15726, W10731);
not G17118 (W15721, W16368);
nor G17119 (W15722, W16369, W16370, W16371);
nor G17120 (W15723, W16372, W16373, W16374);
and G17121 (W15724, W16375, W16376, W16377);
and G17122 (W15725, W16378, W16379, W16380);
and G17123 (W15726, W8185, W16381, I1514);
nor G17124 (W15727, W15728, W13200);
nand G17125 (W15728, W15729, I370);
nor G17126 (W15729, W15730, W13206);
nand G17127 (W15730, W15731, I372);
nor G17128 (W15731, W15732, W13212);
nand G17129 (W15732, W15733, I374);
nor G17130 (W15733, W15734, W13218);
nand G17131 (W15734, W15735, I376);
nor G17132 (W15735, W15736, W13224);
nand G17133 (W15736, W8185, W13640);
not G17134 (W15737, W16382);
not G17135 (W15738, I1515);
not G17136 (W15739, W16383);
not G17137 (W15740, W16384);
not G17138 (W15741, W16385);
not G17139 (W15742, W16386);
nand G17140 (W15743, W16387, W16388);
nand G17141 (W15744, W8243, W16388);
not G17142 (W15745, W16389);
nor G17143 (W15746, W15813, W16390, W14842);
not G17144 (W15747, I1516);
not G17145 (W15748, I157);
not G17146 (W15749, I158);
nor G17147 (W15750, W14840, W16390, W13363);
not G17148 (W15751, W16391);
not G17149 (W15752, I1463);
not G17150 (W15753, W16392);
not G17151 (W15754, I1517);
not G17152 (W15755, W16393);
not G17153 (W15756, W16394);
not G17154 (W15757, W16395);
not G17155 (W15758, W16396);
not G17156 (W15759, W16397);
not G17157 (W15760, W14853);
nor G17158 (W15761, W16398, W16399, W16400);
nor G17159 (W15762, W16401, W16402);
not G17160 (W15763, W16403);
not G17161 (W15764, W16404);
nor G17162 (W15765, W16405, W16406);
not G17163 (W15766, W15768);
nand G17164 (W15767, W11332, W16407);
not G17165 (W15768, W16408);
not G17166 (W15769, I197);
not G17167 (W15770, I196);
nor G17168 (W15771, W16409, W16410);
not G17169 (W15772, W15774);
nor G17170 (W15773, W16411, W16412);
not G17171 (W15774, W16413);
nor G17172 (W15775, W16414, W16415);
not G17173 (W15776, W15778);
nor G17174 (W15777, W16416, W16417);
not G17175 (W15778, W16418);
nor G17176 (W15779, W16419, W16420);
not G17177 (W15780, W15782);
nor G17178 (W15781, W16421, W16422);
not G17179 (W15782, W16423);
nor G17180 (W15783, W16424, W16425);
not G17181 (W15784, W15786);
nand G17182 (W15785, W11328, W16407);
not G17183 (W15786, W16426);
nor G17184 (W15787, W16427, W16428);
not G17185 (W15788, W15790);
nand G17186 (W15789, W11336, W16407);
not G17187 (W15790, W16429);
nor G17188 (W15791, W16430, W16431);
not G17189 (W15792, W15794);
nand G17190 (W15793, W11344, W16407);
not G17191 (W15794, W16432);
nor G17192 (W15795, W16433, W16434);
not G17193 (W15796, W15798);
nor G17194 (W15797, W16435, W16436);
not G17195 (W15798, W16437);
nor G17196 (W15799, W16438, W16439);
not G17197 (W15800, W15802);
nor G17198 (W15801, W16440, W16441);
not G17199 (W15802, W16442);
nor G17200 (W15803, W16443, W16444);
not G17201 (W15804, W15806);
nand G17202 (W15805, W11324, W16407);
not G17203 (W15806, W16445);
nand G17204 (W15807, W16446, W16447);
nand G17205 (W15808, W14842, W16447);
nand G17206 (W15809, W16448, W16449);
nand G17207 (W15810, W16450, W16451);
nand G17208 (W15811, W16390, W16451);
not G17209 (W15812, W16452);
not G17210 (W15813, W16453);
nor G17211 (W15814, W16454, W16455, W16456);
nor G17212 (W15815, W16457, W16458);
not G17213 (W15816, W16459);
not G17214 (W15817, W16460);
nand G17215 (W15818, W16461, W16462, W16463);
not G17216 (W15819, W16453);
not G17217 (W15820, W16464);
not G17218 (W15821, W5386);
nor G17219 (W15822, W14854, W14853);
nor G17220 (W15823, W5394, W5386);
nor G17221 (W15824, W13397, W16465, W13395);
nand G17222 (W15825, W15824, W15751);
and G17223 (W15826, W13417, W11261);
and G17224 (W15827, W13418, W11264);
and G17225 (W15828, W13419, W11267);
not G17226 (W15829, W16466);
not G17227 (W15830, W15751);
not G17228 (W15831, W16467);
or G17229 (W15832, W16468, W11259);
nand G17230 (W15833, W16469, W16470);
nand G17231 (W15834, W15831, W16470);
nor G17232 (W15835, W13395, W16471);
nand G17233 (W15836, W15835, W5385);
nor G17234 (W15837, W13395, W16472);
nand G17235 (W15838, W15837, W15839);
not G17236 (W15839, W16473);
nor G17237 (W15840, W16474, W16475);
not G17238 (W15841, W15839);
not G17239 (W15842, W16476);
or G17240 (W15843, W16477, W14884);
not G17241 (W15844, W16478);
nor G17242 (W15845, W16479, W11428);
nand G17243 (W15846, W15845, I1343);
nor G17244 (W15847, W15846, W13466);
nand G17245 (W15848, W15847, I1345);
nor G17246 (W15849, W15848, W13472);
nand G17247 (W15850, W15849, I1347);
nor G17248 (W15851, W15850, W13478);
nand G17249 (W15852, W15851, I1349);
nor G17250 (W15853, W15852, W13484);
nand G17251 (W15854, W15853, I1351);
not G17252 (W15855, W16480);
not G17253 (W15856, W16481);
not G17254 (W15857, W16482);
not G17255 (W15858, I1518);
not G17256 (W15859, W16483);
not G17257 (W15860, I255);
not G17258 (W15861, W16484);
not G17259 (W15862, W16485);
not G17260 (W15863, W16486);
not G17261 (W15864, W16487);
nand G17262 (W15865, W16488, W16489);
nand G17263 (W15866, W16490, W16489);
nand G17264 (W15867, W16491, W16492);
nand G17265 (W15868, W16493, W16492);
nand G17266 (W15869, W16494, W16495);
nand G17267 (W15870, W16496, W16495);
nand G17268 (W15871, W16497, W16498);
nand G17269 (W15872, W16499, W16498);
and G17270 (W15873, W13569, W13562, I1383, W13559);
and G17271 (W15874, W13587, W13573, W16500);
nand G17272 (W15875, W15877, I1383);
nand G17273 (W15876, W11644, I1384);
nor G17274 (W15877, W15876, W13562);
nor G17275 (W15878, W15883, W13587);
nand G17276 (W15879, W14978, I1391);
nor G17277 (W15880, W15879, W13575);
nand G17278 (W15881, W15880, I1387);
nor G17279 (W15882, W15881, W13581);
nand G17280 (W15883, W15882, I1389);
not G17281 (W15884, W16501);
or G17282 (W15885, W16502, W16503);
or G17283 (W15886, W16504, W16505);
nand G17284 (W15887, W16506, W16507);
nand G17285 (W15888, W15887, W15889);
nand G17286 (W15889, W16508, W16509);
nand G17287 (W15890, W16510, W16511);
nand G17288 (W15891, W15890, W15892);
nand G17289 (W15892, W16512, W16513);
not G17290 (W15893, I1519);
nand G17291 (W15894, W16514, W16515);
nand G17292 (W15895, W15894, W15896);
nand G17293 (W15896, W16516, W16517);
nand G17294 (W15897, W16518, W16519);
nand G17295 (W15898, W15897, W15899);
nand G17296 (W15899, W16520, W16521);
and G17297 (W15900, W11756, W11749, W16522);
and G17298 (W15901, W16523, W16524, W16525);
and G17299 (W15902, W16526, W16527, W16525);
not G17300 (W15903, W13612);
and G17301 (W15904, W16528, W16524, W16529);
and G17302 (W15905, W16526, W16528, W16530);
not G17303 (W15906, W13612);
not G17304 (W15907, W16531);
not G17305 (W15908, I1520);
nor G17306 (W15909, W16532, W16533, W16534);
not G17307 (W15910, I1521);
nor G17308 (W15911, W16535, W16536, W16537);
and G17309 (W15912, W16538, W16539, W16540);
and G17310 (W15913, W16541, W16542, W16540);
not G17311 (W15914, W13619);
and G17312 (W15915, W16543, W16539, W16544);
and G17313 (W15916, W16541, W16543, W16545);
not G17314 (W15917, W13619);
not G17315 (W15918, I1522);
nor G17316 (W15919, W16546, W16547, W16548);
not G17317 (W15920, I1523);
nor G17318 (W15921, W16549, W16550, W16551);
and G17319 (W15922, W16552, W16553, W16554);
and G17320 (W15923, W16555, W16556, W16554);
not G17321 (W15924, W13626);
and G17322 (W15925, W16557, W16553, W16558);
and G17323 (W15926, W16555, W16557, W16559);
not G17324 (W15927, W13626);
not G17325 (W15928, I1524);
nor G17326 (W15929, W16560, W16561, W16562);
not G17327 (W15930, I1525);
nor G17328 (W15931, W16563, W16564, W16565);
and G17329 (W15932, W16566, W16567, W16568);
and G17330 (W15933, W16569, W16570, W16568);
not G17331 (W15934, W13633);
and G17332 (W15935, W16571, W16567, W16572);
and G17333 (W15936, W16569, W16571, W16573);
not G17334 (W15937, W13633);
not G17335 (W15938, I1526);
nor G17336 (W15939, W16574, W16575, W16576);
not G17337 (W15940, I1527);
nor G17338 (W15941, W16577, W16578, W16579);
not G17339 (W15942, W4292);
not G17340 (W15943, W16580);
not G17341 (W15944, W4305);
not G17342 (W15945, W4318);
not G17343 (W15946, W4331);
nand G17344 (W15947, W13783, I1395);
not G17345 (W15948, W16581);
not G17346 (W15949, W16582);
not G17347 (W15950, W15966);
nand G17348 (W15951, W16583, W16584);
not G17349 (W15952, W16585);
not G17350 (W15953, W13815);
not G17351 (W15954, W16586);
not G17352 (W15955, W13815);
nand G17353 (W15956, W16587, W16588);
not G17354 (W15957, W16589);
not G17355 (W15958, W13815);
not G17356 (W15959, W16590);
not G17357 (W15960, W13815);
nand G17358 (W15961, W16591, W16592);
not G17359 (W15962, W16593);
not G17360 (W15963, W13815);
and G17361 (W15964, W16594, W16595);
and G17362 (W15965, W16596, W16597);
nand G17363 (W15966, W16598, W16583);
nand G17364 (W15967, W16599, W16600);
nand G17365 (W15968, W16601, W16600);
nand G17366 (W15969, W16602, W16603);
nand G17367 (W15970, W16604, W16603);
nand G17368 (W15971, W16605, W16606);
not G17369 (W15972, W16607);
not G17370 (W15973, W13815);
not G17371 (W15974, W16608);
not G17372 (W15975, W13815);
not G17373 (W15976, W16609);
not G17374 (W15977, W13815);
not G17375 (W15978, I3);
and G17376 (W15979, W15138, W8440);
and G17377 (W15980, W8544, W8437);
and G17378 (W15981, W13643, W8434);
and G17379 (W15982, W15138, W8450);
and G17380 (W15983, W8544, W8447);
and G17381 (W15984, W13643, W8444);
nand G17382 (W15985, W16610, W16611);
nand G17383 (W15986, W16612, W16613);
and G17384 (W15987, W16614, W16615, W16616);
nand G17385 (W15988, W16617, W16618);
nand G17386 (W15989, W16619, W16620);
and G17387 (W15990, W16621, W16622, W16623);
not G17388 (W15991, W16624);
nor G17389 (W15992, W8372, W16625);
nand G17390 (W15993, W15992, W8372);
not G17391 (W15994, W16062);
nor G17392 (W15995, W16626, W16627, W16628);
and G17393 (W15996, W12210, W8740);
and G17394 (W15997, W12211, W8743);
and G17395 (W15998, W12212, W8746);
or G17396 (W15999, W16629, W16630, W16631);
or G17397 (W16000, W16632, W16633, W16634);
nor G17398 (W16001, W16635, W16636, W16637);
not G17399 (W16002, I1407);
and G17400 (W16003, W16638, W16639);
and G17401 (W16004, W16640, W16641);
or G17402 (W16005, W16642, W16643);
not G17403 (W16006, W16644);
and G17404 (W16007, W16645, W16646);
and G17405 (W16008, W16647, W16648);
and G17406 (W16009, W16649, W16650);
and G17407 (W16010, W9029, W16651);
not G17408 (W16011, W16644);
and G17409 (W16012, W16652, W16653);
and G17410 (W16013, W16654, W16655);
and G17411 (W16014, W16649, W16656);
and G17412 (W16015, W9041, W16657);
not G17413 (W16016, W16644);
and G17414 (W16017, W16658, W16659);
and G17415 (W16018, W16660, W16661);
and G17416 (W16019, W16649, W16662);
and G17417 (W16020, W9009, W16663);
not G17418 (W16021, W16644);
and G17419 (W16022, W16664, W16665);
and G17420 (W16023, W16666, W16667);
not G17421 (W16024, W16644);
and G17422 (W16025, W16668, W16669);
and G17423 (W16026, W16670, W16671);
not G17424 (W16027, W16644);
and G17425 (W16028, W16672, W16673);
and G17426 (W16029, W16674, W16675);
not G17427 (W16030, W16644);
and G17428 (W16031, W16676, W16677);
and G17429 (W16032, W16678, W16679);
and G17430 (W16033, W16649, W16680);
and G17431 (W16034, W9037, W16681);
not G17432 (W16035, W16644);
and G17433 (W16036, W16682, W16683);
and G17434 (W16037, W16684, W16685);
and G17435 (W16038, W16649, W16686);
and G17436 (W16039, W9005, W16687);
not G17437 (W16040, W16644);
and G17438 (W16041, W16688, W16689);
and G17439 (W16042, W16690, W16691);
not G17440 (W16043, W16644);
nor G17441 (W16044, W16692, W16693);
nand G17442 (W16045, W16044, W13984);
nand G17443 (W16046, W16694, W16695);
nand G17444 (W16047, W15244, W16695);
nor G17445 (W16048, W16696, W16697);
nand G17446 (W16049, W16048, W15994);
nand G17447 (W16050, W15193, W15194, W9108, W16698);
nor G17448 (W16051, W16699, W16700, W16701);
and G17449 (W16052, W12210, W8848);
and G17450 (W16053, W12211, W8852);
and G17451 (W16054, W12212, W8855);
and G17452 (W16055, W16702, W16703);
and G17453 (W16056, W12188, W16704);
nor G17454 (W16057, W15244, W15994, W13984);
and G17455 (W16058, W16645, W16678, W16705, W16706);
and G17456 (W16059, W16707, W16708, W16709);
not G17457 (W16060, W12062);
and G17458 (W16061, W16710, W16711, W16712);
nor G17459 (W16062, W16713, W16714, W16715);
not G17460 (W16063, W12189);
nand G17461 (W16064, W16716, W16717);
nor G17462 (W16065, W16718, W16719, W16720);
nor G17463 (W16066, W12188, W16721);
nand G17464 (W16067, W15195, W16722);
nand G17465 (W16068, W16067, W15263);
nor G17466 (W16069, W16723, W16724);
nor G17467 (W16070, W16725, W16726);
nor G17468 (W16071, W16727, W16728, W16729);
and G17469 (W16072, W16730, W16731);
and G17470 (W16073, W16732, W16733);
nor G17471 (W16074, W16734, W16735, W16736);
nor G17472 (W16075, W12188, W15271, W15272);
not G17473 (W16076, W9108);
not G17474 (W16077, I1408);
not G17475 (W16078, W5541);
not G17476 (W16079, W16737);
not G17477 (W16080, W16096);
nand G17478 (W16081, W16738, W16739);
not G17479 (W16082, W16740);
not G17480 (W16083, W14112);
not G17481 (W16084, W16741);
not G17482 (W16085, W14112);
nand G17483 (W16086, W16742, W16743);
not G17484 (W16087, W16744);
not G17485 (W16088, W14112);
not G17486 (W16089, W16745);
not G17487 (W16090, W14112);
nand G17488 (W16091, W16746, W16747);
not G17489 (W16092, W16748);
not G17490 (W16093, W14112);
and G17491 (W16094, W16749, W16750);
and G17492 (W16095, W16751, W16752);
nand G17493 (W16096, W16753, W16738);
nand G17494 (W16097, W16754, W16755);
nand G17495 (W16098, W16756, W16755);
nand G17496 (W16099, W16757, W16758);
nand G17497 (W16100, W16759, W16758);
nand G17498 (W16101, W16760, W16761);
not G17499 (W16102, W16762);
not G17500 (W16103, W14112);
not G17501 (W16104, W16763);
not G17502 (W16105, W14112);
not G17503 (W16106, W16764);
not G17504 (W16107, W14112);
not G17505 (W16108, I52);
and G17506 (W16109, W15335, W9213);
and G17507 (W16110, W9317, W9210);
and G17508 (W16111, W13642, W9207);
and G17509 (W16112, W15335, W9223);
and G17510 (W16113, W9317, W9220);
and G17511 (W16114, W13642, W9217);
nand G17512 (W16115, W16765, W16766);
nand G17513 (W16116, W16767, W16768);
and G17514 (W16117, W16769, W16770, W16771);
nand G17515 (W16118, W16772, W16773);
nand G17516 (W16119, W16774, W16775);
and G17517 (W16120, W16776, W16777, W16778);
not G17518 (W16121, W16779);
nor G17519 (W16122, W8329, W16780);
nand G17520 (W16123, W16122, W8329);
not G17521 (W16124, W16192);
nor G17522 (W16125, W16781, W16782, W16783);
and G17523 (W16126, W12616, W9513);
and G17524 (W16127, W12617, W9516);
and G17525 (W16128, W12618, W9519);
or G17526 (W16129, W16784, W16785, W16786);
or G17527 (W16130, W16787, W16788, W16789);
nor G17528 (W16131, W16790, W16791, W16792);
not G17529 (W16132, I1420);
and G17530 (W16133, W16793, W16794);
and G17531 (W16134, W16795, W16796);
or G17532 (W16135, W16797, W16798);
not G17533 (W16136, W16799);
and G17534 (W16137, W16800, W16801);
and G17535 (W16138, W16802, W16803);
and G17536 (W16139, W16804, W16805);
and G17537 (W16140, W9802, W16806);
not G17538 (W16141, W16799);
and G17539 (W16142, W16807, W16808);
and G17540 (W16143, W16809, W16810);
and G17541 (W16144, W16804, W16811);
and G17542 (W16145, W9814, W16812);
not G17543 (W16146, W16799);
and G17544 (W16147, W16813, W16814);
and G17545 (W16148, W16815, W16816);
and G17546 (W16149, W16804, W16817);
and G17547 (W16150, W9782, W16818);
not G17548 (W16151, W16799);
and G17549 (W16152, W16819, W16820);
and G17550 (W16153, W16821, W16822);
not G17551 (W16154, W16799);
and G17552 (W16155, W16823, W16824);
and G17553 (W16156, W16825, W16826);
not G17554 (W16157, W16799);
and G17555 (W16158, W16827, W16828);
and G17556 (W16159, W16829, W16830);
not G17557 (W16160, W16799);
and G17558 (W16161, W16831, W16832);
and G17559 (W16162, W16833, W16834);
and G17560 (W16163, W16804, W16835);
and G17561 (W16164, W9810, W16836);
not G17562 (W16165, W16799);
and G17563 (W16166, W16837, W16838);
and G17564 (W16167, W16839, W16840);
and G17565 (W16168, W16804, W16841);
and G17566 (W16169, W9778, W16842);
not G17567 (W16170, W16799);
and G17568 (W16171, W16843, W16844);
and G17569 (W16172, W16845, W16846);
not G17570 (W16173, W16799);
nor G17571 (W16174, W16847, W16848);
nand G17572 (W16175, W16174, W14278);
nand G17573 (W16176, W16849, W16850);
nand G17574 (W16177, W15438, W16850);
nor G17575 (W16178, W16851, W16852);
nand G17576 (W16179, W16178, W16124);
nand G17577 (W16180, W15387, W15388, W9881, W16853);
nor G17578 (W16181, W16854, W16855, W16856);
and G17579 (W16182, W12616, W9621);
and G17580 (W16183, W12617, W9625);
and G17581 (W16184, W12618, W9628);
and G17582 (W16185, W16857, W16858);
and G17583 (W16186, W12594, W16859);
nor G17584 (W16187, W15438, W16124, W14278);
and G17585 (W16188, W16800, W16833, W16860, W16861);
and G17586 (W16189, W16862, W16863, W16864);
not G17587 (W16190, W12468);
and G17588 (W16191, W16865, W16866, W16867);
nor G17589 (W16192, W16868, W16869, W16870);
not G17590 (W16193, W12595);
nand G17591 (W16194, W16871, W16872);
nor G17592 (W16195, W16873, W16874, W16875);
nor G17593 (W16196, W12594, W16876);
nand G17594 (W16197, W15389, W16877);
nand G17595 (W16198, W16197, W15456);
nor G17596 (W16199, W16878, W16879);
nor G17597 (W16200, W16880, W16881);
nor G17598 (W16201, W16882, W16883, W16884);
and G17599 (W16202, W16885, W16886);
and G17600 (W16203, W16887, W16888);
nor G17601 (W16204, W16889, W16890, W16891);
nor G17602 (W16205, W12594, W15464, W15465);
not G17603 (W16206, W9881);
not G17604 (W16207, I1421);
not G17605 (W16208, W5540);
not G17606 (W16209, W16892);
not G17607 (W16210, W16226);
nand G17608 (W16211, W16893, W16894);
not G17609 (W16212, W16895);
not G17610 (W16213, W14405);
not G17611 (W16214, W16896);
not G17612 (W16215, W14405);
nand G17613 (W16216, W16897, W16898);
not G17614 (W16217, W16899);
not G17615 (W16218, W14405);
not G17616 (W16219, W16900);
not G17617 (W16220, W14405);
nand G17618 (W16221, W16901, W16902);
not G17619 (W16222, W16903);
not G17620 (W16223, W14405);
and G17621 (W16224, W16904, W16905);
and G17622 (W16225, W16906, W16907);
nand G17623 (W16226, W16908, W16893);
nand G17624 (W16227, W16909, W16910);
nand G17625 (W16228, W16911, W16910);
nand G17626 (W16229, W16912, W16913);
nand G17627 (W16230, W16914, W16913);
nand G17628 (W16231, W16915, W16916);
not G17629 (W16232, W16917);
not G17630 (W16233, W14405);
not G17631 (W16234, W16918);
not G17632 (W16235, W14405);
not G17633 (W16236, W16919);
not G17634 (W16237, W14405);
not G17635 (W16238, I101);
and G17636 (W16239, W15528, W9986);
and G17637 (W16240, W10090, W9983);
and G17638 (W16241, W13641, W9980);
and G17639 (W16242, W15528, W9996);
and G17640 (W16243, W10090, W9993);
and G17641 (W16244, W13641, W9990);
nand G17642 (W16245, W16920, W16921);
nand G17643 (W16246, W16922, W16923);
and G17644 (W16247, W16924, W16925, W16926);
nand G17645 (W16248, W16927, W16928);
nand G17646 (W16249, W16929, W16930);
and G17647 (W16250, W16931, W16932, W16933);
not G17648 (W16251, W16934);
nor G17649 (W16252, W8286, W16935);
nand G17650 (W16253, W16252, W8286);
not G17651 (W16254, W16322);
nor G17652 (W16255, W16936, W16937, W16938);
and G17653 (W16256, W13022, W10286);
and G17654 (W16257, W13023, W10289);
and G17655 (W16258, W13024, W10292);
or G17656 (W16259, W16939, W16940, W16941);
or G17657 (W16260, W16942, W16943, W16944);
nor G17658 (W16261, W16945, W16946, W16947);
not G17659 (W16262, I1433);
and G17660 (W16263, W16948, W16949);
and G17661 (W16264, W16950, W16951);
or G17662 (W16265, W16952, W16953);
not G17663 (W16266, W16954);
and G17664 (W16267, W16955, W16956);
and G17665 (W16268, W16957, W16958);
and G17666 (W16269, W16959, W16960);
and G17667 (W16270, W10571, W16961);
not G17668 (W16271, W16954);
and G17669 (W16272, W16962, W16963);
and G17670 (W16273, W16964, W16965);
and G17671 (W16274, W16959, W16966);
and G17672 (W16275, W10583, W16967);
not G17673 (W16276, W16954);
and G17674 (W16277, W16968, W16969);
and G17675 (W16278, W16970, W16971);
and G17676 (W16279, W16959, W16972);
and G17677 (W16280, W10551, W16973);
not G17678 (W16281, W16954);
and G17679 (W16282, W16974, W16975);
and G17680 (W16283, W16976, W16977);
not G17681 (W16284, W16954);
and G17682 (W16285, W16978, W16979);
and G17683 (W16286, W16980, W16981);
not G17684 (W16287, W16954);
and G17685 (W16288, W16982, W16983);
and G17686 (W16289, W16984, W16985);
not G17687 (W16290, W16954);
and G17688 (W16291, W16986, W16987);
and G17689 (W16292, W16988, W16989);
and G17690 (W16293, W16959, W16990);
and G17691 (W16294, W10579, W16991);
not G17692 (W16295, W16954);
and G17693 (W16296, W16992, W16993);
and G17694 (W16297, W16994, W16995);
and G17695 (W16298, W16959, W16996);
and G17696 (W16299, W10587, W16997);
not G17697 (W16300, W16954);
and G17698 (W16301, W16998, W16999);
and G17699 (W16302, W17000, W17001);
not G17700 (W16303, W16954);
nor G17701 (W16304, W17002, W17003);
nand G17702 (W16305, W16304, W14571);
nand G17703 (W16306, W17004, W17005);
nand G17704 (W16307, W15631, W17005);
nor G17705 (W16308, W17006, W17007);
nand G17706 (W16309, W16308, W16254);
nand G17707 (W16310, W15580, W15581, W10654, W17008);
nor G17708 (W16311, W17009, W17010, W17011);
and G17709 (W16312, W13022, W10394);
and G17710 (W16313, W13023, W10398);
and G17711 (W16314, W13024, W10401);
and G17712 (W16315, W17012, W17013);
and G17713 (W16316, W13000, W17014);
nor G17714 (W16317, W15631, W16254, W14571);
and G17715 (W16318, W16955, W16988, W17015, W17016);
and G17716 (W16319, W17017, W17018, W17019);
not G17717 (W16320, W12874);
and G17718 (W16321, W17020, W17021, W17022);
nor G17719 (W16322, W17023, W17024, W17025);
not G17720 (W16323, W13001);
nand G17721 (W16324, W17026, W17027);
nor G17722 (W16325, W17028, W17029, W17030);
nor G17723 (W16326, W13000, W17031);
nand G17724 (W16327, W15582, W17032);
nand G17725 (W16328, W16327, W15649);
nor G17726 (W16329, W17033, W17034);
nor G17727 (W16330, W17035, W17036);
nor G17728 (W16331, W17037, W17038, W17039);
and G17729 (W16332, W17040, W17041);
and G17730 (W16333, W17042, W17043);
nor G17731 (W16334, W17044, W17045, W17046);
nor G17732 (W16335, W13000, W15657, W15658);
not G17733 (W16336, W10654);
not G17734 (W16337, I1434);
not G17735 (W16338, W5539);
not G17736 (W16339, W17047);
not G17737 (W16340, W16356);
nand G17738 (W16341, W17048, W17049);
not G17739 (W16342, W17050);
not G17740 (W16343, W14698);
not G17741 (W16344, W17051);
not G17742 (W16345, W14698);
nand G17743 (W16346, W17052, W17053);
not G17744 (W16347, W17054);
not G17745 (W16348, W14698);
not G17746 (W16349, W17055);
not G17747 (W16350, W14698);
nand G17748 (W16351, W17056, W17057);
not G17749 (W16352, W17058);
not G17750 (W16353, W14698);
and G17751 (W16354, W17059, W17060);
and G17752 (W16355, W17061, W17062);
nand G17753 (W16356, W17063, W17048);
nand G17754 (W16357, W17064, W17065);
nand G17755 (W16358, W17066, W17065);
nand G17756 (W16359, W17067, W17068);
nand G17757 (W16360, W17069, W17068);
nand G17758 (W16361, W17070, W17071);
not G17759 (W16362, W17072);
not G17760 (W16363, W14698);
not G17761 (W16364, W17073);
not G17762 (W16365, W14698);
not G17763 (W16366, W17074);
not G17764 (W16367, W14698);
not G17765 (W16368, I150);
and G17766 (W16369, W15721, W10759);
and G17767 (W16370, W10863, W10756);
and G17768 (W16371, W13640, W10753);
and G17769 (W16372, W15721, W10769);
and G17770 (W16373, W10863, W10766);
and G17771 (W16374, W13640, W10763);
nand G17772 (W16375, W17075, W17076);
nand G17773 (W16376, W17077, W17078);
and G17774 (W16377, W17079, W17080, W17081);
nand G17775 (W16378, W17082, W17083);
nand G17776 (W16379, W17084, W17085);
and G17777 (W16380, W17086, W17087, W17088);
not G17778 (W16381, W17089);
not G17779 (W16382, W11016);
not G17780 (W16383, W11016);
not G17781 (W16384, W11016);
not G17782 (W16385, W11016);
not G17783 (W16386, W11016);
nor G17784 (W16387, W8243, W17090);
nand G17785 (W16388, W16387, W8243);
not G17786 (W16389, W11015);
not G17787 (W16390, W16464);
nor G17788 (W16391, W17091, W17092, W17093);
not G17789 (W16392, W13418);
not G17790 (W16393, W13418);
not G17791 (W16394, W13418);
not G17792 (W16395, W13418);
not G17793 (W16396, W13418);
not G17794 (W16397, W13418);
and G17795 (W16398, W13417, W11059);
and G17796 (W16399, W13418, W11062);
and G17797 (W16400, W13419, W11065);
or G17798 (W16401, W17094, W17095, W17096);
or G17799 (W16402, W17097, W17098, W17099);
nor G17800 (W16403, W17100, W17101, W17102);
not G17801 (W16404, I1446);
and G17802 (W16405, W17103, W17104);
and G17803 (W16406, W17105, W17106);
or G17804 (W16407, W17107, W17108);
not G17805 (W16408, W17109);
and G17806 (W16409, W17110, W17111);
and G17807 (W16410, W17112, W17113);
and G17808 (W16411, W17114, W17115);
and G17809 (W16412, W11340, W17116);
not G17810 (W16413, W17109);
and G17811 (W16414, W17117, W17118);
and G17812 (W16415, W17119, W17120);
and G17813 (W16416, W17114, W17121);
and G17814 (W16417, W11352, W17122);
not G17815 (W16418, W17109);
and G17816 (W16419, W17123, W17124);
and G17817 (W16420, W17125, W17126);
and G17818 (W16421, W17114, W17127);
and G17819 (W16422, W11363, W17128);
not G17820 (W16423, W17109);
and G17821 (W16424, W17129, W17130);
and G17822 (W16425, W17131, W17132);
not G17823 (W16426, W17109);
and G17824 (W16427, W17133, W17134);
and G17825 (W16428, W17135, W17136);
not G17826 (W16429, W17109);
and G17827 (W16430, W17137, W17138);
and G17828 (W16431, W17139, W17140);
not G17829 (W16432, W17109);
and G17830 (W16433, W17141, W17142);
and G17831 (W16434, W17143, W17144);
and G17832 (W16435, W17114, W17145);
and G17833 (W16436, W11348, W17146);
not G17834 (W16437, W17109);
and G17835 (W16438, W17147, W17148);
and G17836 (W16439, W17149, W17150);
and G17837 (W16440, W17114, W17151);
and G17838 (W16441, W11356, W17152);
not G17839 (W16442, W17109);
and G17840 (W16443, W17153, W17154);
and G17841 (W16444, W17155, W17156);
not G17842 (W16445, W17109);
nor G17843 (W16446, W17157, W17158);
nand G17844 (W16447, W16446, W14842);
nand G17845 (W16448, W17159, W17160);
nand G17846 (W16449, W15813, W17160);
nor G17847 (W16450, W17161, W17162);
nand G17848 (W16451, W16450, W16390);
nand G17849 (W16452, W15762, W15763, W11427, W17163);
nor G17850 (W16453, W17164, W17165, W17166);
and G17851 (W16454, W13417, W11167);
and G17852 (W16455, W13418, W11171);
and G17853 (W16456, W13419, W11174);
and G17854 (W16457, W17167, W17168);
and G17855 (W16458, W13395, W17169);
nor G17856 (W16459, W15813, W16390, W14842);
and G17857 (W16460, W17110, W17143, W17170, W17171);
and G17858 (W16461, W17172, W17173, W17174);
not G17859 (W16462, W13275);
and G17860 (W16463, W17175, W17176, W17177);
nor G17861 (W16464, W17178, W17179, W17180);
not G17862 (W16465, W13396);
nand G17863 (W16466, W17181, W17182);
nor G17864 (W16467, W17183, W17184, W17185);
nor G17865 (W16468, W13395, W17186);
nand G17866 (W16469, W15764, W17187);
nand G17867 (W16470, W16469, W15831);
nor G17868 (W16471, W17188, W17189);
nor G17869 (W16472, W17190, W17191);
nor G17870 (W16473, W17192, W17193, W17194);
and G17871 (W16474, W17195, W17196);
and G17872 (W16475, W17197, W17198);
nor G17873 (W16476, W17199, W17200, W17201);
nor G17874 (W16477, W13395, W15839, W15840);
not G17875 (W16478, W11427);
not G17876 (W16479, I1447);
not G17877 (W16480, W5538);
or G17878 (W16481, W17202, W17203);
or G17879 (W16482, W17204, W17205);
not G17880 (W16483, I255);
or G17881 (W16484, W17206, W17207);
or G17882 (W16485, W17208, W17209);
or G17883 (W16486, W17210, W17211);
or G17884 (W16487, W17212, W17213);
nand G17885 (W16488, W17214, W17215);
nand G17886 (W16489, W16488, W16490);
nand G17887 (W16490, W17216, W17217);
nand G17888 (W16491, W17218, W17219);
nand G17889 (W16492, W16491, W16493);
nand G17890 (W16493, W17220, W17221);
nand G17891 (W16494, W17222, W17223);
nand G17892 (W16495, W16494, W16496);
nand G17893 (W16496, W17224, W17225);
nand G17894 (W16497, W17226, W17227);
nand G17895 (W16498, W16497, W16499);
nand G17896 (W16499, W17228, W17229);
and G17897 (W16500, W13579, W13581, W13585);
not G17898 (W16501, I1528);
and G17899 (W16502, W17230, W17231);
not G17900 (W16503, W17230);
and G17901 (W16504, W17230, W17232);
not G17902 (W16505, W17230);
nand G17903 (W16506, W17233, W17234);
nand G17904 (W16507, W17235, W17234);
nand G17905 (W16508, W17236, W17237);
nand G17906 (W16509, W17238, W17237);
nand G17907 (W16510, W17239, W17240);
nand G17908 (W16511, W17241, W17240);
nand G17909 (W16512, W17242, W17243);
nand G17910 (W16513, W17244, W17243);
nand G17911 (W16514, W17245, W17246);
nand G17912 (W16515, W17247, W17246);
nand G17913 (W16516, W17248, W17249);
nand G17914 (W16517, W17250, W17249);
nand G17915 (W16518, W17251, W17252);
nand G17916 (W16519, W17253, W17252);
nand G17917 (W16520, W17254, W17255);
nand G17918 (W16521, W17256, W17255);
and G17919 (W16522, W13782, I503, I501);
not G17920 (W16523, W16526);
nor G17921 (W16524, W15005, W15004);
not G17922 (W16525, W16529);
nor G17923 (W16526, W15003, W15002);
or G17924 (W16527, W17257, W17258);
not G17925 (W16528, W16527);
or G17926 (W16529, W17259, W17260, W17261);
not G17927 (W16530, W16524);
not G17928 (W16531, W17262);
and G17929 (W16532, W11015, I458);
and G17930 (W16533, W11016, I459);
and G17931 (W16534, W11017, I460);
and G17932 (W16535, W11015, I461);
and G17933 (W16536, W11016, I462);
and G17934 (W16537, W11017, I463);
not G17935 (W16538, W16541);
nor G17936 (W16539, W15018, W15017);
not G17937 (W16540, W16544);
nor G17938 (W16541, W15016, W15015);
or G17939 (W16542, W17263, W17264);
not G17940 (W16543, W16542);
or G17941 (W16544, W17265, W17266, W17267);
not G17942 (W16545, W16539);
and G17943 (W16546, W10242, I470);
and G17944 (W16547, W10243, I471);
and G17945 (W16548, W10244, I472);
and G17946 (W16549, W10242, I473);
and G17947 (W16550, W10243, I474);
and G17948 (W16551, W10244, I475);
not G17949 (W16552, W16555);
nor G17950 (W16553, W15031, W15030);
not G17951 (W16554, W16558);
nor G17952 (W16555, W15029, W15028);
or G17953 (W16556, W17268, W17269);
not G17954 (W16557, W16556);
or G17955 (W16558, W17270, W17271, W17272);
not G17956 (W16559, W16553);
and G17957 (W16560, W9469, I482);
and G17958 (W16561, W9470, I483);
and G17959 (W16562, W9471, I484);
and G17960 (W16563, W9469, I485);
and G17961 (W16564, W9470, I486);
and G17962 (W16565, W9471, I487);
not G17963 (W16566, W16569);
nor G17964 (W16567, W15044, W15043);
not G17965 (W16568, W16572);
nor G17966 (W16569, W15042, W15041);
or G17967 (W16570, W17273, W17274);
not G17968 (W16571, W16570);
or G17969 (W16572, W17275, W17276, W17277);
not G17970 (W16573, W16567);
and G17971 (W16574, W8696, I494);
and G17972 (W16575, W8697, I495);
and G17973 (W16576, W8698, I496);
and G17974 (W16577, W8696, I497);
and G17975 (W16578, W8697, I498);
and G17976 (W16579, W8698, I499);
not G17977 (W16580, W17278);
not G17978 (W16581, I1529);
or G17979 (W16582, W17279, I1449, W4435);
nand G17980 (W16583, W17280, W17281, W17282);
nand G17981 (W16584, W11867, W17282);
nand G17982 (W16585, W17283, W17284);
nand G17983 (W16586, W17285, W17286);
not G17984 (W16587, W17287);
not G17985 (W16588, W17288);
nand G17986 (W16589, W17289, W17290);
nand G17987 (W16590, W17291, W17292);
nand G17988 (W16591, W8432, W17293);
nand G17989 (W16592, W17294, W17293);
nand G17990 (W16593, W17295, W17296);
not G17991 (W16594, I1477);
not G17992 (W16595, W16597);
not G17993 (W16596, I1530);
not G17994 (W16597, W17297);
nand G17995 (W16598, W11917, W17281);
nand G17996 (W16599, W17298, W17299);
nand G17997 (W16600, W16599, W16601);
nand G17998 (W16601, W17300, W17301);
nand G17999 (W16602, W17302, W17303);
nand G18000 (W16603, W16602, W16604);
nand G18001 (W16604, W17304, W17305);
nand G18002 (W16605, W8442, W17306);
nand G18003 (W16606, W17307, W17306);
nand G18004 (W16607, W17308, W17309);
nand G18005 (W16608, W17310, W17311);
nand G18006 (W16609, W17312, W17313);
nand G18007 (W16610, W11982, W17314);
nand G18008 (W16611, W17315, W17314);
nand G18009 (W16612, W11979, W17316);
nand G18010 (W16613, W17317, W17316);
nand G18011 (W16614, W17318, W17319);
nand G18012 (W16615, W17320, W17321);
nand G18013 (W16616, W17322, W17323);
nand G18014 (W16617, W11998, W17324);
nand G18015 (W16618, W17325, W17324);
nand G18016 (W16619, W11994, W17326);
nand G18017 (W16620, W17327, W17326);
nand G18018 (W16621, W17328, W17329);
nand G18019 (W16622, W17330, W17331);
nand G18020 (W16623, W17332, W17333);
not G18021 (W16624, I1531);
and G18022 (W16625, W17334, W11867);
and G18023 (W16626, W12210, I692);
and G18024 (W16627, W12211, I693);
and G18025 (W16628, W12212, I694);
nand G18026 (W16629, W17335, W17336);
nand G18027 (W16630, W17337, W17338);
or G18028 (W16631, W17339, W17340, W17341);
nand G18029 (W16632, W17342, W17343);
nand G18030 (W16633, W17344, W17345);
or G18031 (W16634, W17346, W17347, W17348);
and G18032 (W16635, W13950, W9164);
and G18033 (W16636, W13951, W9161);
and G18034 (W16637, W9107, W9158);
not G18035 (W16638, W16640);
not G18036 (W16639, W16641);
not G18037 (W16640, W17349);
not G18038 (W16641, W17350);
not G18039 (W16642, W17351);
nand G18040 (W16643, W17352, W17353);
or G18041 (W16644, W16643, W17351);
not G18042 (W16645, W16647);
not G18043 (W16646, W16648);
not G18044 (W16647, W17354);
not G18045 (W16648, W17355);
not G18046 (W16649, W17356);
not G18047 (W16650, W16651);
not G18048 (W16651, W17357);
not G18049 (W16652, W16654);
not G18050 (W16653, W16655);
not G18051 (W16654, W17358);
not G18052 (W16655, W17359);
not G18053 (W16656, W16657);
not G18054 (W16657, W17360);
not G18055 (W16658, W17361);
not G18056 (W16659, W16661);
not G18057 (W16660, W16658);
not G18058 (W16661, W17362);
not G18059 (W16662, W16663);
not G18060 (W16663, W17363);
not G18061 (W16664, W17364);
not G18062 (W16665, W16667);
not G18063 (W16666, W16664);
not G18064 (W16667, W17365);
not G18065 (W16668, W17366);
not G18066 (W16669, W16671);
not G18067 (W16670, W16668);
not G18068 (W16671, W17367);
not G18069 (W16672, W17368);
not G18070 (W16673, W16675);
not G18071 (W16674, W16672);
not G18072 (W16675, W17369);
not G18073 (W16676, W17370);
not G18074 (W16677, W16679);
not G18075 (W16678, W16676);
not G18076 (W16679, W17371);
not G18077 (W16680, W16681);
not G18078 (W16681, W17372);
not G18079 (W16682, W16684);
not G18080 (W16683, W16685);
not G18081 (W16684, W17373);
not G18082 (W16685, W17374);
not G18083 (W16686, W16687);
not G18084 (W16687, W17375);
not G18085 (W16688, W16690);
not G18086 (W16689, W16691);
not G18087 (W16690, W17376);
not G18088 (W16691, W17377);
and G18089 (W16692, W17378, W17379);
and G18090 (W16693, W17380, W17381);
nor G18091 (W16694, W17382, W17383);
nand G18092 (W16695, W16694, W15244);
and G18093 (W16696, W17384, W17385);
and G18094 (W16697, W17386, W17387);
and G18095 (W16698, W17388, W17389);
and G18096 (W16699, W12210, W8858);
and G18097 (W16700, W12211, W8862);
and G18098 (W16701, W12212, W8865);
not G18099 (W16702, W17390);
not G18100 (W16703, W16704);
not G18101 (W16704, W17391);
and G18102 (W16705, W16638, W16670, W17392);
and G18103 (W16706, W16652, W16682, W16660);
nand G18104 (W16707, W17393, W17394);
nand G18105 (W16708, W17395, W17396);
and G18106 (W16709, W17397, W17398, W17399);
nand G18107 (W16710, W17400, W17401);
nand G18108 (W16711, W17402, W17403);
and G18109 (W16712, W17404, W17405, W17406);
and G18110 (W16713, W12210, W8868);
and G18111 (W16714, W12211, W8872);
and G18112 (W16715, W12212, W8875);
not G18113 (W16716, W17407);
and G18114 (W16717, W17408, W17409);
and G18115 (W16718, W12210, I699);
and G18116 (W16719, W12211, I700);
and G18117 (W16720, W12212, I698);
nor G18118 (W16721, W17410, W17411);
nand G18119 (W16722, W17412, W17413);
and G18120 (W16723, W17414, W17415);
and G18121 (W16724, W17416, W17417);
and G18122 (W16725, W17418, W17419);
and G18123 (W16726, W17420, W17421);
and G18124 (W16727, W12210, I704);
and G18125 (W16728, W12211, I705);
and G18126 (W16729, W12212, I706);
nor G18127 (W16730, W16732, W17422);
not G18128 (W16731, W16733);
not G18129 (W16732, W17423);
not G18130 (W16733, W17424);
and G18131 (W16734, W12210, W8982);
and G18132 (W16735, W12211, W8985);
and G18133 (W16736, W12212, W8988);
or G18134 (W16737, W17425, I1453, W4710);
nand G18135 (W16738, W17426, W17427, W17428);
nand G18136 (W16739, W11841, W17428);
nand G18137 (W16740, W17429, W17430);
nand G18138 (W16741, W17431, W17432);
not G18139 (W16742, W17433);
not G18140 (W16743, W17434);
nand G18141 (W16744, W17435, W17436);
nand G18142 (W16745, W17437, W17438);
nand G18143 (W16746, W9205, W17439);
nand G18144 (W16747, W17440, W17439);
nand G18145 (W16748, W17441, W17442);
not G18146 (W16749, I1490);
not G18147 (W16750, W16752);
not G18148 (W16751, I1532);
not G18149 (W16752, W17443);
nand G18150 (W16753, W12323, W17427);
nand G18151 (W16754, W17444, W17445);
nand G18152 (W16755, W16754, W16756);
nand G18153 (W16756, W17446, W17447);
nand G18154 (W16757, W17448, W17449);
nand G18155 (W16758, W16757, W16759);
nand G18156 (W16759, W17450, W17451);
nand G18157 (W16760, W9215, W17452);
nand G18158 (W16761, W17453, W17452);
nand G18159 (W16762, W17454, W17455);
nand G18160 (W16763, W17456, W17457);
nand G18161 (W16764, W17458, W17459);
nand G18162 (W16765, W12388, W17460);
nand G18163 (W16766, W17461, W17460);
nand G18164 (W16767, W12385, W17462);
nand G18165 (W16768, W17463, W17462);
nand G18166 (W16769, W17464, W17465);
nand G18167 (W16770, W17466, W17467);
nand G18168 (W16771, W17468, W17469);
nand G18169 (W16772, W12404, W17470);
nand G18170 (W16773, W17471, W17470);
nand G18171 (W16774, W12400, W17472);
nand G18172 (W16775, W17473, W17472);
nand G18173 (W16776, W17474, W17475);
nand G18174 (W16777, W17476, W17477);
nand G18175 (W16778, W17478, W17479);
not G18176 (W16779, I1533);
and G18177 (W16780, W17480, W11841);
and G18178 (W16781, W12616, I893);
and G18179 (W16782, W12617, I894);
and G18180 (W16783, W12618, I895);
nand G18181 (W16784, W17481, W17482);
nand G18182 (W16785, W17483, W17484);
or G18183 (W16786, W17485, W17486, W17487);
nand G18184 (W16787, W17488, W17489);
nand G18185 (W16788, W17490, W17491);
or G18186 (W16789, W17492, W17493, W17494);
and G18187 (W16790, W14244, W9937);
and G18188 (W16791, W14245, W9934);
and G18189 (W16792, W9880, W9931);
not G18190 (W16793, W16795);
not G18191 (W16794, W16796);
not G18192 (W16795, W17495);
not G18193 (W16796, W17496);
not G18194 (W16797, W17497);
nand G18195 (W16798, W17498, W17499);
or G18196 (W16799, W16798, W17497);
not G18197 (W16800, W16802);
not G18198 (W16801, W16803);
not G18199 (W16802, W17500);
not G18200 (W16803, W17501);
not G18201 (W16804, W17502);
not G18202 (W16805, W16806);
not G18203 (W16806, W17503);
not G18204 (W16807, W16809);
not G18205 (W16808, W16810);
not G18206 (W16809, W17504);
not G18207 (W16810, W17505);
not G18208 (W16811, W16812);
not G18209 (W16812, W17506);
not G18210 (W16813, W17507);
not G18211 (W16814, W16816);
not G18212 (W16815, W16813);
not G18213 (W16816, W17508);
not G18214 (W16817, W16818);
not G18215 (W16818, W17509);
not G18216 (W16819, W17510);
not G18217 (W16820, W16822);
not G18218 (W16821, W16819);
not G18219 (W16822, W17511);
not G18220 (W16823, W17512);
not G18221 (W16824, W16826);
not G18222 (W16825, W16823);
not G18223 (W16826, W17513);
not G18224 (W16827, W17514);
not G18225 (W16828, W16830);
not G18226 (W16829, W16827);
not G18227 (W16830, W17515);
not G18228 (W16831, W17516);
not G18229 (W16832, W16834);
not G18230 (W16833, W16831);
not G18231 (W16834, W17517);
not G18232 (W16835, W16836);
not G18233 (W16836, W17518);
not G18234 (W16837, W16839);
not G18235 (W16838, W16840);
not G18236 (W16839, W17519);
not G18237 (W16840, W17520);
not G18238 (W16841, W16842);
not G18239 (W16842, W17521);
not G18240 (W16843, W16845);
not G18241 (W16844, W16846);
not G18242 (W16845, W17522);
not G18243 (W16846, W17523);
and G18244 (W16847, W17524, W17525);
and G18245 (W16848, W17526, W17527);
nor G18246 (W16849, W17528, W17529);
nand G18247 (W16850, W16849, W15438);
and G18248 (W16851, W17530, W17531);
and G18249 (W16852, W17532, W17533);
and G18250 (W16853, W17534, W17535);
and G18251 (W16854, W12616, W9631);
and G18252 (W16855, W12617, W9635);
and G18253 (W16856, W12618, W9638);
not G18254 (W16857, W17536);
not G18255 (W16858, W16859);
not G18256 (W16859, W17537);
and G18257 (W16860, W16793, W16825, W17538);
and G18258 (W16861, W16807, W16837, W16815);
nand G18259 (W16862, W17539, W17540);
nand G18260 (W16863, W17541, W17542);
and G18261 (W16864, W17543, W17544, W17545);
nand G18262 (W16865, W17546, W17547);
nand G18263 (W16866, W17548, W17549);
and G18264 (W16867, W17550, W17551, W17552);
and G18265 (W16868, W12616, W9641);
and G18266 (W16869, W12617, W9645);
and G18267 (W16870, W12618, W9648);
not G18268 (W16871, W17553);
and G18269 (W16872, W17554, W17555);
and G18270 (W16873, W12616, I900);
and G18271 (W16874, W12617, I901);
and G18272 (W16875, W12618, I899);
nor G18273 (W16876, W17556, W17557);
nand G18274 (W16877, W17558, W17559);
and G18275 (W16878, W17560, W17561);
and G18276 (W16879, W17562, W17563);
and G18277 (W16880, W17564, W17565);
and G18278 (W16881, W17566, W17567);
and G18279 (W16882, W12616, I905);
and G18280 (W16883, W12617, I906);
and G18281 (W16884, W12618, I907);
nor G18282 (W16885, W16887, W17568);
not G18283 (W16886, W16888);
not G18284 (W16887, W17569);
not G18285 (W16888, W17570);
and G18286 (W16889, W12616, W9755);
and G18287 (W16890, W12617, W9758);
and G18288 (W16891, W12618, W9761);
or G18289 (W16892, W17571, I1457, W4985);
nand G18290 (W16893, W17572, W17573, W17574);
nand G18291 (W16894, W11815, W17574);
nand G18292 (W16895, W17575, W17576);
nand G18293 (W16896, W17577, W17578);
not G18294 (W16897, W17579);
not G18295 (W16898, W17580);
nand G18296 (W16899, W17581, W17582);
nand G18297 (W16900, W17583, W17584);
nand G18298 (W16901, W9978, W17585);
nand G18299 (W16902, W17586, W17585);
nand G18300 (W16903, W17587, W17588);
not G18301 (W16904, I1502);
not G18302 (W16905, W16907);
not G18303 (W16906, I1534);
not G18304 (W16907, W17589);
nand G18305 (W16908, W12729, W17573);
nand G18306 (W16909, W17590, W17591);
nand G18307 (W16910, W16909, W16911);
nand G18308 (W16911, W17592, W17593);
nand G18309 (W16912, W17594, W17595);
nand G18310 (W16913, W16912, W16914);
nand G18311 (W16914, W17596, W17597);
nand G18312 (W16915, W9988, W17598);
nand G18313 (W16916, W17599, W17598);
nand G18314 (W16917, W17600, W17601);
nand G18315 (W16918, W17602, W17603);
nand G18316 (W16919, W17604, W17605);
nand G18317 (W16920, W12794, W17606);
nand G18318 (W16921, W17607, W17606);
nand G18319 (W16922, W12791, W17608);
nand G18320 (W16923, W17609, W17608);
nand G18321 (W16924, W17610, W17611);
nand G18322 (W16925, W17612, W17613);
nand G18323 (W16926, W17614, W17615);
nand G18324 (W16927, W12810, W17616);
nand G18325 (W16928, W17617, W17616);
nand G18326 (W16929, W12806, W17618);
nand G18327 (W16930, W17619, W17618);
nand G18328 (W16931, W17620, W17621);
nand G18329 (W16932, W17622, W17623);
nand G18330 (W16933, W17624, W17625);
not G18331 (W16934, I1535);
and G18332 (W16935, W17626, W11815);
and G18333 (W16936, W13022, I1094);
and G18334 (W16937, W13023, I1095);
and G18335 (W16938, W13024, I1096);
nand G18336 (W16939, W17627, W17628);
nand G18337 (W16940, W17629, W17630);
or G18338 (W16941, W17631, W17632, W17633);
nand G18339 (W16942, W17634, W17635);
nand G18340 (W16943, W17636, W17637);
or G18341 (W16944, W17638, W17639, W17640);
and G18342 (W16945, W14537, W10710);
and G18343 (W16946, W14538, W10707);
and G18344 (W16947, W10653, W10704);
not G18345 (W16948, W16950);
not G18346 (W16949, W16951);
not G18347 (W16950, W17641);
not G18348 (W16951, W17642);
not G18349 (W16952, W17643);
nand G18350 (W16953, W17644, W17645);
or G18351 (W16954, W16953, W17643);
not G18352 (W16955, W16957);
not G18353 (W16956, W16958);
not G18354 (W16957, W17646);
not G18355 (W16958, W17647);
not G18356 (W16959, W17648);
not G18357 (W16960, W16961);
not G18358 (W16961, W17649);
not G18359 (W16962, W16964);
not G18360 (W16963, W16965);
not G18361 (W16964, W17650);
not G18362 (W16965, W17651);
not G18363 (W16966, W16967);
not G18364 (W16967, W17652);
not G18365 (W16968, W17653);
not G18366 (W16969, W16971);
not G18367 (W16970, W16968);
not G18368 (W16971, W17654);
not G18369 (W16972, W16973);
not G18370 (W16973, W17655);
not G18371 (W16974, W17656);
not G18372 (W16975, W16977);
not G18373 (W16976, W16974);
not G18374 (W16977, W17657);
not G18375 (W16978, W17658);
not G18376 (W16979, W16981);
not G18377 (W16980, W16978);
not G18378 (W16981, W17659);
not G18379 (W16982, W17660);
not G18380 (W16983, W16985);
not G18381 (W16984, W16982);
not G18382 (W16985, W17661);
not G18383 (W16986, W17662);
not G18384 (W16987, W16989);
not G18385 (W16988, W16986);
not G18386 (W16989, W17663);
not G18387 (W16990, W16991);
not G18388 (W16991, W17664);
not G18389 (W16992, W16994);
not G18390 (W16993, W16995);
not G18391 (W16994, W17665);
not G18392 (W16995, W17666);
not G18393 (W16996, W16997);
not G18394 (W16997, W17667);
not G18395 (W16998, W17000);
not G18396 (W16999, W17001);
not G18397 (W17000, W17668);
not G18398 (W17001, W17669);
and G18399 (W17002, W17670, W17671);
and G18400 (W17003, W17672, W17673);
nor G18401 (W17004, W17674, W17675);
nand G18402 (W17005, W17004, W15631);
and G18403 (W17006, W17676, W17677);
and G18404 (W17007, W17678, W17679);
and G18405 (W17008, W17680, W17681);
and G18406 (W17009, W13022, W10404);
and G18407 (W17010, W13023, W10408);
and G18408 (W17011, W13024, W10411);
not G18409 (W17012, W17682);
not G18410 (W17013, W17014);
not G18411 (W17014, W17683);
and G18412 (W17015, W16948, W16980, W17684);
and G18413 (W17016, W16962, W16992, W16970);
nand G18414 (W17017, W17685, W17686);
nand G18415 (W17018, W17687, W17688);
and G18416 (W17019, W17689, W17690, W17691);
nand G18417 (W17020, W17692, W17693);
nand G18418 (W17021, W17694, W17695);
and G18419 (W17022, W17696, W17697, W17698);
and G18420 (W17023, W13022, W10414);
and G18421 (W17024, W13023, W10418);
and G18422 (W17025, W13024, W10421);
not G18423 (W17026, W17699);
and G18424 (W17027, W17700, W17701);
and G18425 (W17028, W13022, I1101);
and G18426 (W17029, W13023, I1102);
and G18427 (W17030, W13024, I1100);
nor G18428 (W17031, W17702, W17703);
nand G18429 (W17032, W17704, W17705);
and G18430 (W17033, W17706, W17707);
and G18431 (W17034, W17708, W17709);
and G18432 (W17035, W17710, W17711);
and G18433 (W17036, W17712, W17713);
and G18434 (W17037, W13022, I1106);
and G18435 (W17038, W13023, I1107);
and G18436 (W17039, W13024, I1108);
nor G18437 (W17040, W17042, W17714);
not G18438 (W17041, W17043);
not G18439 (W17042, W17715);
not G18440 (W17043, W17716);
and G18441 (W17044, W13022, W10528);
and G18442 (W17045, W13023, W10531);
and G18443 (W17046, W13024, W10534);
or G18444 (W17047, W17717, I1461, W17718, W5260);
nand G18445 (W17048, W17719, W17720, W17721);
nand G18446 (W17049, W11788, W17721);
nand G18447 (W17050, W17722, W17723);
nand G18448 (W17051, W17724, W17725);
not G18449 (W17052, W17726);
not G18450 (W17053, W17727);
nand G18451 (W17054, W17728, W17729);
nand G18452 (W17055, W17730, W17731);
nand G18453 (W17056, W10751, W17732);
nand G18454 (W17057, W17733, W17732);
nand G18455 (W17058, W17734, W17735);
not G18456 (W17059, I1514);
not G18457 (W17060, W17062);
not G18458 (W17061, I1536);
not G18459 (W17062, W17736);
nand G18460 (W17063, W13135, W17720);
nand G18461 (W17064, W17737, W17738);
nand G18462 (W17065, W17064, W17066);
nand G18463 (W17066, W17739, W17740);
nand G18464 (W17067, W17741, W17742);
nand G18465 (W17068, W17067, W17069);
nand G18466 (W17069, W17743, W17744);
nand G18467 (W17070, W10761, W17745);
nand G18468 (W17071, W17746, W17745);
nand G18469 (W17072, W17747, W17748);
nand G18470 (W17073, W17749, W17750);
nand G18471 (W17074, W17751, W17752);
nand G18472 (W17075, W13200, W17753);
nand G18473 (W17076, W17754, W17753);
nand G18474 (W17077, W13197, W17755);
nand G18475 (W17078, W17756, W17755);
nand G18476 (W17079, W17757, W17758);
nand G18477 (W17080, W17759, W17760);
nand G18478 (W17081, W17761, W17762);
nand G18479 (W17082, W13216, W17763);
nand G18480 (W17083, W17764, W17763);
nand G18481 (W17084, W13212, W17765);
nand G18482 (W17085, W17766, W17765);
nand G18483 (W17086, W17767, W17768);
nand G18484 (W17087, W17769, W17770);
nand G18485 (W17088, W17771, W17772);
not G18486 (W17089, I1537);
and G18487 (W17090, W17773, W11788);
and G18488 (W17091, W13417, I1295);
and G18489 (W17092, W13418, I1296);
and G18490 (W17093, W13419, I1297);
nand G18491 (W17094, W17774, W17775);
nand G18492 (W17095, W17776, W17777);
or G18493 (W17096, W17778, W17779, W17780);
nand G18494 (W17097, W17781, W17782);
nand G18495 (W17098, W17783, W17784);
or G18496 (W17099, W17785, W17786, W17787);
and G18497 (W17100, W14808, W11483);
and G18498 (W17101, W14809, W11480);
and G18499 (W17102, W11426, W11477);
not G18500 (W17103, W17105);
not G18501 (W17104, W17106);
not G18502 (W17105, W17788);
not G18503 (W17106, W17789);
not G18504 (W17107, W17790);
nand G18505 (W17108, W17791, W17792);
or G18506 (W17109, W17108, W17790);
not G18507 (W17110, W17112);
not G18508 (W17111, W17113);
not G18509 (W17112, W17793);
not G18510 (W17113, W17794);
not G18511 (W17114, W17795);
not G18512 (W17115, W17116);
not G18513 (W17116, W17796);
not G18514 (W17117, W17119);
not G18515 (W17118, W17120);
not G18516 (W17119, W17797);
not G18517 (W17120, W17798);
not G18518 (W17121, W17122);
not G18519 (W17122, W17799);
not G18520 (W17123, W17800);
not G18521 (W17124, W17126);
not G18522 (W17125, W17123);
not G18523 (W17126, W17801);
not G18524 (W17127, W17128);
not G18525 (W17128, W17802);
not G18526 (W17129, W17803);
not G18527 (W17130, W17132);
not G18528 (W17131, W17129);
not G18529 (W17132, W17804);
not G18530 (W17133, W17805);
not G18531 (W17134, W17136);
not G18532 (W17135, W17133);
not G18533 (W17136, W17806);
not G18534 (W17137, W17807);
not G18535 (W17138, W17140);
not G18536 (W17139, W17137);
not G18537 (W17140, W17808);
not G18538 (W17141, W17809);
not G18539 (W17142, W17144);
not G18540 (W17143, W17141);
not G18541 (W17144, W17810);
not G18542 (W17145, W17146);
not G18543 (W17146, W17811);
not G18544 (W17147, W17149);
not G18545 (W17148, W17150);
not G18546 (W17149, W17812);
not G18547 (W17150, W17813);
not G18548 (W17151, W17152);
not G18549 (W17152, W17814);
not G18550 (W17153, W17155);
not G18551 (W17154, W17156);
not G18552 (W17155, W17815);
not G18553 (W17156, W17816);
and G18554 (W17157, W17817, W17818);
and G18555 (W17158, W17819, W17820);
nor G18556 (W17159, W17821, W17822);
nand G18557 (W17160, W17159, W15813);
and G18558 (W17161, W17823, W17824);
and G18559 (W17162, W17825, W17826);
and G18560 (W17163, W17827, W17828);
and G18561 (W17164, W13417, W11177);
and G18562 (W17165, W13418, W11181);
and G18563 (W17166, W13419, W11184);
not G18564 (W17167, W17829);
not G18565 (W17168, W17169);
not G18566 (W17169, W17830);
and G18567 (W17170, W17103, W17135, W17831);
and G18568 (W17171, W17117, W17147, W17125);
nand G18569 (W17172, W17832, W17833);
nand G18570 (W17173, W17834, W17835);
and G18571 (W17174, W17836, W17837, W17838);
nand G18572 (W17175, W17839, W17840);
nand G18573 (W17176, W17841, W17842);
and G18574 (W17177, W17843, W17844, W17845);
and G18575 (W17178, W13417, W11187);
and G18576 (W17179, W13418, W11191);
and G18577 (W17180, W13419, W11194);
not G18578 (W17181, W17846);
and G18579 (W17182, W17847, W17848);
and G18580 (W17183, W13417, I1302);
and G18581 (W17184, W13418, I1303);
and G18582 (W17185, W13419, I1301);
nor G18583 (W17186, W17849, W17850);
nand G18584 (W17187, W17851, W17852);
and G18585 (W17188, W17853, W17854);
and G18586 (W17189, W17855, W17856);
and G18587 (W17190, W17857, W17858);
and G18588 (W17191, W17859, W17860);
and G18589 (W17192, W13417, I1307);
and G18590 (W17193, W13418, I1308);
and G18591 (W17194, W13419, I1309);
nor G18592 (W17195, W17197, W17861);
not G18593 (W17196, W17198);
not G18594 (W17197, W17862);
not G18595 (W17198, W17863);
and G18596 (W17199, W13417, W11301);
and G18597 (W17200, W13418, W11304);
and G18598 (W17201, W13419, W11307);
and G18599 (W17202, W17230, W17864);
not G18600 (W17203, W17230);
and G18601 (W17204, W17230, W17865);
not G18602 (W17205, W17230);
and G18603 (W17206, W17230, W17866);
not G18604 (W17207, W17230);
and G18605 (W17208, W17230, W17867);
not G18606 (W17209, W17230);
and G18607 (W17210, W17230, W17868);
not G18608 (W17211, W17230);
and G18609 (W17212, W17230, W17869);
not G18610 (W17213, W17230);
nand G18611 (W17214, I1365, W17870);
nand G18612 (W17215, I1366, W17870);
nand G18613 (W17216, I1367, W17871);
nand G18614 (W17217, I1368, W17871);
nand G18615 (W17218, I1369, W17872);
nand G18616 (W17219, I1370, W17872);
nand G18617 (W17220, I1371, W17873);
nand G18618 (W17221, I1372, W17873);
nand G18619 (W17222, I1373, W17874);
nand G18620 (W17223, I1374, W17874);
nand G18621 (W17224, I1375, W17875);
nand G18622 (W17225, I1376, W17875);
nand G18623 (W17226, I1377, W17876);
nand G18624 (W17227, I1378, W17876);
nand G18625 (W17228, I1379, W17877);
nand G18626 (W17229, I1380, W17877);
not G18627 (W17230, W17878);
not G18628 (W17231, W17879);
not G18629 (W17232, W17880);
not G18630 (W17233, I1538);
nand G18631 (W17234, W17233, W17235);
not G18632 (W17235, I1539);
not G18633 (W17236, I1540);
nand G18634 (W17237, W17236, W17238);
not G18635 (W17238, I1541);
not G18636 (W17239, I1542);
nand G18637 (W17240, W17239, W17241);
not G18638 (W17241, I1543);
not G18639 (W17242, I1544);
nand G18640 (W17243, W17242, W17244);
not G18641 (W17244, I1545);
not G18642 (W17245, I1546);
nand G18643 (W17246, W17245, W17247);
not G18644 (W17247, I1547);
not G18645 (W17248, I1548);
nand G18646 (W17249, W17248, W17250);
not G18647 (W17250, I1549);
not G18648 (W17251, I1550);
nand G18649 (W17252, W17251, W17253);
not G18650 (W17253, I1551);
not G18651 (W17254, I1552);
nand G18652 (W17255, W17254, W17256);
not G18653 (W17256, I1553);
or G18654 (W17257, W17881, W17882, W17883, W17884);
or G18655 (W17258, W17885, W17886, W17887, W17888);
or G18656 (W17259, W17889, W17890, W17891, W17892);
or G18657 (W17260, W17893, W17894, W17895);
or G18658 (W17261, W17896, W17897, W17898);
not G18659 (W17262, I1554);
or G18660 (W17263, W17899, W17900, W17901, W17902);
or G18661 (W17264, W17903, W17904, W17905, W17906);
or G18662 (W17265, W17907, W17908, W17909, W17910);
or G18663 (W17266, W17911, W17912, W17913);
or G18664 (W17267, W17914, W17915, W17916);
or G18665 (W17268, W17917, W17918, W17919, W17920);
or G18666 (W17269, W17921, W17922, W17923, W17924);
or G18667 (W17270, W17925, W17926, W17927, W17928);
or G18668 (W17271, W17929, W17930, W17931);
or G18669 (W17272, W17932, W17933, W17934);
or G18670 (W17273, W17935, W17936, W17937, W17938);
or G18671 (W17274, W17939, W17940, W17941, W17942);
or G18672 (W17275, W17943, W17944, W17945, W17946);
or G18673 (W17276, W17947, W17948, W17949);
or G18674 (W17277, W17950, W17951, W17952);
not G18675 (W17278, W17953);
not G18676 (W17279, W17954);
not G18677 (W17280, W17955);
not G18678 (W17281, W11867);
not G18679 (W17282, W11917);
nand G18680 (W17283, W8442, W17956);
nand G18681 (W17284, W17957, W17956);
nand G18682 (W17285, W8432, W17958);
nand G18683 (W17286, W17959, W17958);
not G18684 (W17287, W17960);
not G18685 (W17288, W17961);
nand G18686 (W17289, W8432, W17962);
nand G18687 (W17290, W17963, W17962);
nand G18688 (W17291, W8442, W17964);
nand G18689 (W17292, W17965, W17964);
nand G18690 (W17293, W8432, W17294);
nand G18691 (W17294, W16588, W17317);
nand G18692 (W17295, W8432, W17966);
nand G18693 (W17296, W17967, W17966);
not G18694 (W17297, W13756);
nand G18695 (W17298, W15125, W17968);
nand G18696 (W17299, W15113, W17968);
nand G18697 (W17300, W15133, W17969);
nand G18698 (W17301, W15129, W17969);
nand G18699 (W17302, W15107, W17970);
nand G18700 (W17303, W15098, W17970);
nand G18701 (W17304, W15094, W17971);
nand G18702 (W17305, W15103, W17971);
nand G18703 (W17306, W8442, W17307);
nand G18704 (W17307, W16588, W17315);
nand G18705 (W17308, W8442, W17972);
nand G18706 (W17309, W17973, W17972);
nand G18707 (W17310, W8432, W17974);
nand G18708 (W17311, W17975, W17974);
nand G18709 (W17312, W8442, W17976);
nand G18710 (W17313, W17977, W17976);
nand G18711 (W17314, W11982, W17315);
not G18712 (W17315, W17978);
nand G18713 (W17316, W11979, W17317);
not G18714 (W17317, W17979);
nand G18715 (W17318, W11992, W17980);
nand G18716 (W17319, W17981, W17980);
nand G18717 (W17320, W11988, W17982);
nand G18718 (W17321, W17983, W17982);
nand G18719 (W17322, W11986, W17984);
nand G18720 (W17323, W17985, W17984);
nand G18721 (W17324, W11998, W17325);
not G18722 (W17325, W17986);
nand G18723 (W17326, W11994, W17327);
not G18724 (W17327, W17987);
nand G18725 (W17328, W12006, W17988);
nand G18726 (W17329, W17989, W17988);
nand G18727 (W17330, W12004, W17990);
nand G18728 (W17331, W17991, W17990);
nand G18729 (W17332, W12000, W17992);
nand G18730 (W17333, W17993, W17992);
not G18731 (W17334, W11866);
nand G18732 (W17335, W9009, W17994);
nand G18733 (W17336, W17995, W17994);
nand G18734 (W17337, W9013, W17996);
nand G18735 (W17338, W17997, W17996);
nand G18736 (W17339, W17998, W17999);
nand G18737 (W17340, W18000, W18001);
nand G18738 (W17341, W18002, W18003);
nand G18739 (W17342, W9029, W18004);
nand G18740 (W17343, W18005, W18004);
nand G18741 (W17344, W9037, W18006);
nand G18742 (W17345, W18007, W18006);
nand G18743 (W17346, W18008, W18009);
nand G18744 (W17347, W18010, W18011);
nand G18745 (W17348, W18012, W18013);
nor G18746 (W17349, W18014, W18015, W18016);
not G18747 (W17350, W18017);
nor G18748 (W17351, W18018, W18019);
not G18749 (W17352, W13970);
nor G18750 (W17353, W18020, W18021, W18022);
nor G18751 (W17354, W18023, W18024, W18025);
not G18752 (W17355, W18026);
not G18753 (W17356, W18027);
not G18754 (W17357, W16005);
nor G18755 (W17358, W18028, W18029, W18030);
not G18756 (W17359, W18031);
not G18757 (W17360, W16005);
nor G18758 (W17361, W18032, W18033, W18034);
not G18759 (W17362, W18035);
not G18760 (W17363, W16005);
nor G18761 (W17364, W18036, W18037, W18038);
not G18762 (W17365, W18039);
nor G18763 (W17366, W18040, W18041, W18042);
not G18764 (W17367, W18043);
nor G18765 (W17368, W18044, W18045, W18046);
not G18766 (W17369, W18047);
nor G18767 (W17370, W18048, W18049, W18050);
not G18768 (W17371, W18051);
not G18769 (W17372, W16005);
nor G18770 (W17373, W18052, W18053, W18054);
not G18771 (W17374, W18055);
not G18772 (W17375, W16005);
nor G18773 (W17376, W18056, W18057, W18058);
not G18774 (W17377, W18059);
nand G18775 (W17378, W18060, W18061);
not G18776 (W17379, W17381);
nor G18777 (W17380, W15244, W13983);
not G18778 (W17381, W18062);
and G18779 (W17382, W18063, W18064);
and G18780 (W17383, W13982, W18065);
nor G18781 (W17384, W18066, W18067);
not G18782 (W17385, W17387);
nand G18783 (W17386, W13983, W13982);
not G18784 (W17387, W18068);
nand G18785 (W17388, W18069, W15194, W9108);
nand G18786 (W17389, W18070, W15194, W9108);
not G18787 (W17390, W18071);
not G18788 (W17391, W15175);
and G18789 (W17392, W16674, W16688, W16666);
nand G18790 (W17393, I743, W18072);
nand G18791 (W17394, W16660, W18072);
nand G18792 (W17395, I744, W18073);
nand G18793 (W17396, W16688, W18073);
nand G18794 (W17397, W18074, W18075);
nand G18795 (W17398, W18076, W18077);
nand G18796 (W17399, W18078, W18079);
nand G18797 (W17400, I748, W18080);
nand G18798 (W17401, W16645, W18080);
nand G18799 (W17402, I749, W18081);
nand G18800 (W17403, W16678, W18081);
nand G18801 (W17404, W18082, W18083);
nand G18802 (W17405, W18084, W18085);
nand G18803 (W17406, W18086, W18087);
nor G18804 (W17407, W18088, W18089, W18090);
and G18805 (W17408, W18091, W18092, W18093, W18094);
and G18806 (W17409, W18095, W18096, W18097, W18098);
nor G18807 (W17410, W18099, W15263, W15176);
and G18808 (W17411, W18099, W15263, W15176);
nand G18809 (W17412, W15263, W18100);
nand G18810 (W17413, W15261, W18100);
nor G18811 (W17414, W18101, W18102);
not G18812 (W17415, W17417);
nor G18813 (W17416, W18103, W18104);
not G18814 (W17417, W18105);
nor G18815 (W17418, W18106, W18107);
not G18816 (W17419, W17421);
nor G18817 (W17420, W18108, W18109);
not G18818 (W17421, W18110);
not G18819 (W17422, W18111);
not G18820 (W17423, W18112);
not G18821 (W17424, W4560);
not G18822 (W17425, W18113);
not G18823 (W17426, W18114);
not G18824 (W17427, W11841);
not G18825 (W17428, W12323);
nand G18826 (W17429, W9215, W18115);
nand G18827 (W17430, W18116, W18115);
nand G18828 (W17431, W9205, W18117);
nand G18829 (W17432, W18118, W18117);
not G18830 (W17433, W18119);
not G18831 (W17434, W18120);
nand G18832 (W17435, W9205, W18121);
nand G18833 (W17436, W18122, W18121);
nand G18834 (W17437, W9215, W18123);
nand G18835 (W17438, W18124, W18123);
nand G18836 (W17439, W9205, W17440);
nand G18837 (W17440, W16743, W17463);
nand G18838 (W17441, W9205, W18125);
nand G18839 (W17442, W18126, W18125);
not G18840 (W17443, W13722);
nand G18841 (W17444, W15322, W18127);
nand G18842 (W17445, W15310, W18127);
nand G18843 (W17446, W15330, W18128);
nand G18844 (W17447, W15326, W18128);
nand G18845 (W17448, W15304, W18129);
nand G18846 (W17449, W15295, W18129);
nand G18847 (W17450, W15291, W18130);
nand G18848 (W17451, W15300, W18130);
nand G18849 (W17452, W9215, W17453);
nand G18850 (W17453, W16743, W17461);
nand G18851 (W17454, W9215, W18131);
nand G18852 (W17455, W18132, W18131);
nand G18853 (W17456, W9205, W18133);
nand G18854 (W17457, W18134, W18133);
nand G18855 (W17458, W9215, W18135);
nand G18856 (W17459, W18136, W18135);
nand G18857 (W17460, W12388, W17461);
not G18858 (W17461, W18137);
nand G18859 (W17462, W12385, W17463);
not G18860 (W17463, W18138);
nand G18861 (W17464, W12398, W18139);
nand G18862 (W17465, W18140, W18139);
nand G18863 (W17466, W12394, W18141);
nand G18864 (W17467, W18142, W18141);
nand G18865 (W17468, W12392, W18143);
nand G18866 (W17469, W18144, W18143);
nand G18867 (W17470, W12404, W17471);
not G18868 (W17471, W18145);
nand G18869 (W17472, W12400, W17473);
not G18870 (W17473, W18146);
nand G18871 (W17474, W12412, W18147);
nand G18872 (W17475, W18148, W18147);
nand G18873 (W17476, W12410, W18149);
nand G18874 (W17477, W18150, W18149);
nand G18875 (W17478, W12406, W18151);
nand G18876 (W17479, W18152, W18151);
not G18877 (W17480, W11840);
nand G18878 (W17481, W9782, W18153);
nand G18879 (W17482, W18154, W18153);
nand G18880 (W17483, W9786, W18155);
nand G18881 (W17484, W18156, W18155);
nand G18882 (W17485, W18157, W18158);
nand G18883 (W17486, W18159, W18160);
nand G18884 (W17487, W18161, W18162);
nand G18885 (W17488, W9802, W18163);
nand G18886 (W17489, W18164, W18163);
nand G18887 (W17490, W9810, W18165);
nand G18888 (W17491, W18166, W18165);
nand G18889 (W17492, W18167, W18168);
nand G18890 (W17493, W18169, W18170);
nand G18891 (W17494, W18171, W18172);
nor G18892 (W17495, W18173, W18174, W18175);
not G18893 (W17496, W18176);
nor G18894 (W17497, W18177, W18178);
not G18895 (W17498, W14264);
nor G18896 (W17499, W18179, W18180, W18181);
nor G18897 (W17500, W18182, W18183, W18184);
not G18898 (W17501, W18185);
not G18899 (W17502, W18186);
not G18900 (W17503, W16135);
nor G18901 (W17504, W18187, W18188, W18189);
not G18902 (W17505, W18190);
not G18903 (W17506, W16135);
nor G18904 (W17507, W18191, W18192, W18193);
not G18905 (W17508, W18194);
not G18906 (W17509, W16135);
nor G18907 (W17510, W18195, W18196, W18197);
not G18908 (W17511, W18198);
nor G18909 (W17512, W18199, W18200, W18201);
not G18910 (W17513, W18202);
nor G18911 (W17514, W18203, W18204, W18205);
not G18912 (W17515, W18206);
nor G18913 (W17516, W18207, W18208, W18209);
not G18914 (W17517, W18210);
not G18915 (W17518, W16135);
nor G18916 (W17519, W18211, W18212, W18213);
not G18917 (W17520, W18214);
not G18918 (W17521, W16135);
nor G18919 (W17522, W18215, W18216, W18217);
not G18920 (W17523, W18218);
nand G18921 (W17524, W18219, W18220);
not G18922 (W17525, W17527);
nor G18923 (W17526, W15438, W14277);
not G18924 (W17527, W18221);
and G18925 (W17528, W18222, W18223);
and G18926 (W17529, W14276, W18224);
nor G18927 (W17530, W18225, W18226);
not G18928 (W17531, W17533);
nand G18929 (W17532, W14277, W14276);
not G18930 (W17533, W18227);
nand G18931 (W17534, W18228, W15388, W9881);
nand G18932 (W17535, W18229, W15388, W9881);
not G18933 (W17536, W18230);
not G18934 (W17537, W15369);
and G18935 (W17538, W16829, W16843, W16821);
nand G18936 (W17539, I944, W18231);
nand G18937 (W17540, W16815, W18231);
nand G18938 (W17541, I945, W18232);
nand G18939 (W17542, W16843, W18232);
nand G18940 (W17543, W18233, W18234);
nand G18941 (W17544, W18235, W18236);
nand G18942 (W17545, W18237, W18238);
nand G18943 (W17546, I949, W18239);
nand G18944 (W17547, W16800, W18239);
nand G18945 (W17548, I950, W18240);
nand G18946 (W17549, W16833, W18240);
nand G18947 (W17550, W18241, W18242);
nand G18948 (W17551, W18243, W18244);
nand G18949 (W17552, W18245, W18246);
nor G18950 (W17553, W18247, W18248, W18249);
and G18951 (W17554, W18250, W18251, W18252, W18253);
and G18952 (W17555, W18254, W18255, W18256, W18257);
nor G18953 (W17556, W18258, W15456, W15370);
and G18954 (W17557, W18258, W15456, W15370);
nand G18955 (W17558, W15456, W18259);
nand G18956 (W17559, W15454, W18259);
nor G18957 (W17560, W18260, W18261);
not G18958 (W17561, W17563);
nor G18959 (W17562, W18262, W18263);
not G18960 (W17563, W18264);
nor G18961 (W17564, W18265, W18266);
not G18962 (W17565, W17567);
nor G18963 (W17566, W18267, W18268);
not G18964 (W17567, W18269);
not G18965 (W17568, W18270);
not G18966 (W17569, W18271);
not G18967 (W17570, W4835);
not G18968 (W17571, W18272);
not G18969 (W17572, W18273);
not G18970 (W17573, W11815);
not G18971 (W17574, W12729);
nand G18972 (W17575, W9988, W18274);
nand G18973 (W17576, W18275, W18274);
nand G18974 (W17577, W9978, W18276);
nand G18975 (W17578, W18277, W18276);
not G18976 (W17579, W18278);
not G18977 (W17580, W18279);
nand G18978 (W17581, W9978, W18280);
nand G18979 (W17582, W18281, W18280);
nand G18980 (W17583, W9988, W18282);
nand G18981 (W17584, W18283, W18282);
nand G18982 (W17585, W9978, W17586);
nand G18983 (W17586, W16898, W17609);
nand G18984 (W17587, W9978, W18284);
nand G18985 (W17588, W18285, W18284);
not G18986 (W17589, W13688);
nand G18987 (W17590, W15515, W18286);
nand G18988 (W17591, W15503, W18286);
nand G18989 (W17592, W15523, W18287);
nand G18990 (W17593, W15519, W18287);
nand G18991 (W17594, W15497, W18288);
nand G18992 (W17595, W15488, W18288);
nand G18993 (W17596, W15484, W18289);
nand G18994 (W17597, W15493, W18289);
nand G18995 (W17598, W9988, W17599);
nand G18996 (W17599, W16898, W17607);
nand G18997 (W17600, W9988, W18290);
nand G18998 (W17601, W18291, W18290);
nand G18999 (W17602, W9978, W18292);
nand G19000 (W17603, W18293, W18292);
nand G19001 (W17604, W9988, W18294);
nand G19002 (W17605, W18295, W18294);
nand G19003 (W17606, W12794, W17607);
not G19004 (W17607, W18296);
nand G19005 (W17608, W12791, W17609);
not G19006 (W17609, W18297);
nand G19007 (W17610, W12804, W18298);
nand G19008 (W17611, W18299, W18298);
nand G19009 (W17612, W12800, W18300);
nand G19010 (W17613, W18301, W18300);
nand G19011 (W17614, W12798, W18302);
nand G19012 (W17615, W18303, W18302);
nand G19013 (W17616, W12810, W17617);
not G19014 (W17617, W18304);
nand G19015 (W17618, W12806, W17619);
not G19016 (W17619, W18305);
nand G19017 (W17620, W12818, W18306);
nand G19018 (W17621, W18307, W18306);
nand G19019 (W17622, W12816, W18308);
nand G19020 (W17623, W18309, W18308);
nand G19021 (W17624, W12812, W18310);
nand G19022 (W17625, W18311, W18310);
not G19023 (W17626, W11814);
nand G19024 (W17627, W10551, W18312);
nand G19025 (W17628, W18313, W18312);
nand G19026 (W17629, W10555, W18314);
nand G19027 (W17630, W18315, W18314);
nand G19028 (W17631, W18316, W18317);
nand G19029 (W17632, W18318, W18319);
nand G19030 (W17633, W18320, W18321);
nand G19031 (W17634, W10571, W18322);
nand G19032 (W17635, W18323, W18322);
nand G19033 (W17636, W10579, W18324);
nand G19034 (W17637, W18325, W18324);
nand G19035 (W17638, W18326, W18327);
nand G19036 (W17639, W18328, W18329);
nand G19037 (W17640, W18330, W18331);
nor G19038 (W17641, W18332, W18333, W18334);
not G19039 (W17642, W18335);
nor G19040 (W17643, W18336, W18337);
not G19041 (W17644, W14557);
nor G19042 (W17645, W18338, W18339, W18340);
nor G19043 (W17646, W18341, W18342, W18343);
not G19044 (W17647, W18344);
not G19045 (W17648, W18345);
not G19046 (W17649, W16265);
nor G19047 (W17650, W18346, W18347, W18348);
not G19048 (W17651, W18349);
not G19049 (W17652, W16265);
nor G19050 (W17653, W18350, W18351, W18352);
not G19051 (W17654, W18353);
not G19052 (W17655, W16265);
nor G19053 (W17656, W18354, W18355, W18356);
not G19054 (W17657, W18357);
nor G19055 (W17658, W18358, W18359, W18360);
not G19056 (W17659, W18361);
nor G19057 (W17660, W18362, W18363, W18364);
not G19058 (W17661, W18365);
nor G19059 (W17662, W18366, W18367, W18368);
not G19060 (W17663, W18369);
not G19061 (W17664, W16265);
nor G19062 (W17665, W18370, W18371, W18372);
not G19063 (W17666, W18373);
not G19064 (W17667, W16265);
nor G19065 (W17668, W18374, W18375, W18376);
not G19066 (W17669, W18377);
nand G19067 (W17670, W18378, W18379);
not G19068 (W17671, W17673);
nor G19069 (W17672, W15631, W14570);
not G19070 (W17673, W18380);
and G19071 (W17674, W18381, W18382);
and G19072 (W17675, W14569, W18383);
nor G19073 (W17676, W18384, W18385);
not G19074 (W17677, W17679);
nand G19075 (W17678, W14570, W14569);
not G19076 (W17679, W18386);
nand G19077 (W17680, W18387, W15581, W10654);
nand G19078 (W17681, W18388, W15581, W10654);
not G19079 (W17682, W18389);
not G19080 (W17683, W15562);
and G19081 (W17684, W16984, W16998, W16976);
nand G19082 (W17685, I1145, W18390);
nand G19083 (W17686, W16970, W18390);
nand G19084 (W17687, I1146, W18391);
nand G19085 (W17688, W16998, W18391);
nand G19086 (W17689, W18392, W18393);
nand G19087 (W17690, W18394, W18395);
nand G19088 (W17691, W18396, W18397);
nand G19089 (W17692, I1150, W18398);
nand G19090 (W17693, W16955, W18398);
nand G19091 (W17694, I1151, W18399);
nand G19092 (W17695, W16988, W18399);
nand G19093 (W17696, W18400, W18401);
nand G19094 (W17697, W18402, W18403);
nand G19095 (W17698, W18404, W18405);
nor G19096 (W17699, W18406, W18407, W18408);
and G19097 (W17700, W18409, W18410, W18411, W18412);
and G19098 (W17701, W18413, W18414, W18415, W18416);
nor G19099 (W17702, W18417, W15649, W15563);
and G19100 (W17703, W18417, W15649, W15563);
nand G19101 (W17704, W15649, W18418);
nand G19102 (W17705, W15647, W18418);
nor G19103 (W17706, W18419, W18420);
not G19104 (W17707, W17709);
nor G19105 (W17708, W18421, W18422);
not G19106 (W17709, W18423);
nor G19107 (W17710, W18424, W18425);
not G19108 (W17711, W17713);
nor G19109 (W17712, W18426, W18427);
not G19110 (W17713, W18428);
not G19111 (W17714, W18429);
not G19112 (W17715, W18430);
not G19113 (W17716, W5110);
not G19114 (W17717, W18431);
nor G19115 (W17718, I222, W18432);
not G19116 (W17719, W18433);
not G19117 (W17720, W11788);
not G19118 (W17721, W13135);
nand G19119 (W17722, W10761, W18434);
nand G19120 (W17723, W18435, W18434);
nand G19121 (W17724, W10751, W18436);
nand G19122 (W17725, W18437, W18436);
not G19123 (W17726, W18438);
not G19124 (W17727, W18439);
nand G19125 (W17728, W10751, W18440);
nand G19126 (W17729, W18441, W18440);
nand G19127 (W17730, W10761, W18442);
nand G19128 (W17731, W18443, W18442);
nand G19129 (W17732, W10751, W17733);
nand G19130 (W17733, W17053, W17756);
nand G19131 (W17734, W10751, W18444);
nand G19132 (W17735, W18445, W18444);
not G19133 (W17736, W13653);
nand G19134 (W17737, W15708, W18446);
nand G19135 (W17738, W15696, W18446);
nand G19136 (W17739, W15716, W18447);
nand G19137 (W17740, W15712, W18447);
nand G19138 (W17741, W15690, W18448);
nand G19139 (W17742, W15681, W18448);
nand G19140 (W17743, W15677, W18449);
nand G19141 (W17744, W15686, W18449);
nand G19142 (W17745, W10761, W17746);
nand G19143 (W17746, W17053, W17754);
nand G19144 (W17747, W10761, W18450);
nand G19145 (W17748, W18451, W18450);
nand G19146 (W17749, W10751, W18452);
nand G19147 (W17750, W18453, W18452);
nand G19148 (W17751, W10761, W18454);
nand G19149 (W17752, W18455, W18454);
nand G19150 (W17753, W13200, W17754);
not G19151 (W17754, W18456);
nand G19152 (W17755, W13197, W17756);
not G19153 (W17756, W18457);
nand G19154 (W17757, W13210, W18458);
nand G19155 (W17758, W18459, W18458);
nand G19156 (W17759, W13206, W18460);
nand G19157 (W17760, W18461, W18460);
nand G19158 (W17761, W13204, W18462);
nand G19159 (W17762, W18463, W18462);
nand G19160 (W17763, W13216, W17764);
not G19161 (W17764, W18464);
nand G19162 (W17765, W13212, W17766);
not G19163 (W17766, W18465);
nand G19164 (W17767, W13224, W18466);
nand G19165 (W17768, W18467, W18466);
nand G19166 (W17769, W13222, W18468);
nand G19167 (W17770, W18469, W18468);
nand G19168 (W17771, W13218, W18470);
nand G19169 (W17772, W18471, W18470);
not G19170 (W17773, W11787);
nand G19171 (W17774, W11363, W18472);
nand G19172 (W17775, W18473, W18472);
nand G19173 (W17776, W11324, W18474);
nand G19174 (W17777, W18475, W18474);
nand G19175 (W17778, W18476, W18477);
nand G19176 (W17779, W18478, W18479);
nand G19177 (W17780, W18480, W18481);
nand G19178 (W17781, W11340, W18482);
nand G19179 (W17782, W18483, W18482);
nand G19180 (W17783, W11348, W18484);
nand G19181 (W17784, W18485, W18484);
nand G19182 (W17785, W18486, W18487);
nand G19183 (W17786, W18488, W18489);
nand G19184 (W17787, W18490, W18491);
nor G19185 (W17788, W18492, W18493, W18494);
not G19186 (W17789, W18495);
nor G19187 (W17790, W18496, W18497);
not G19188 (W17791, W14828);
nor G19189 (W17792, W18498, W18499, W18500);
nor G19190 (W17793, W18501, W18502, W18503);
not G19191 (W17794, W18504);
not G19192 (W17795, W18505);
not G19193 (W17796, W16407);
nor G19194 (W17797, W18506, W18507, W18508);
not G19195 (W17798, W18509);
not G19196 (W17799, W16407);
nor G19197 (W17800, W18510, W18511, W18512);
not G19198 (W17801, W18513);
not G19199 (W17802, W16407);
nor G19200 (W17803, W18514, W18515, W18516);
not G19201 (W17804, W18517);
nor G19202 (W17805, W18518, W18519, W18520);
not G19203 (W17806, W18521);
nor G19204 (W17807, W18522, W18523, W18524);
not G19205 (W17808, W18525);
nor G19206 (W17809, W18526, W18527, W18528);
not G19207 (W17810, W18529);
not G19208 (W17811, W16407);
nor G19209 (W17812, W18530, W18531, W18532);
not G19210 (W17813, W18533);
not G19211 (W17814, W16407);
nor G19212 (W17815, W18534, W18535, W18536);
not G19213 (W17816, W18537);
nand G19214 (W17817, W18538, W18539);
not G19215 (W17818, W17820);
nor G19216 (W17819, W15813, W14841);
not G19217 (W17820, W18540);
and G19218 (W17821, W18541, W18542);
and G19219 (W17822, W14840, W18543);
nor G19220 (W17823, W18544, W18545);
not G19221 (W17824, W17826);
nand G19222 (W17825, W14841, W14840);
not G19223 (W17826, W18546);
nand G19224 (W17827, W18547, W15763, W11427);
nand G19225 (W17828, W18548, W15763, W11427);
not G19226 (W17829, W18549);
not G19227 (W17830, W15750);
and G19228 (W17831, W17139, W17153, W17131);
nand G19229 (W17832, I1346, W18550);
nand G19230 (W17833, W17125, W18550);
nand G19231 (W17834, I1347, W18551);
nand G19232 (W17835, W17153, W18551);
nand G19233 (W17836, W18552, W18553);
nand G19234 (W17837, W18554, W18555);
nand G19235 (W17838, W18556, W18557);
nand G19236 (W17839, I1351, W18558);
nand G19237 (W17840, W17110, W18558);
nand G19238 (W17841, I1352, W18559);
nand G19239 (W17842, W17143, W18559);
nand G19240 (W17843, W18560, W18561);
nand G19241 (W17844, W18562, W18563);
nand G19242 (W17845, W18564, W18565);
nor G19243 (W17846, W18566, W18567, W18568);
and G19244 (W17847, W18569, W18570, W18571, W18572);
and G19245 (W17848, W18573, W18574, W18575, W18576);
nor G19246 (W17849, W18577, W15831, W15751);
and G19247 (W17850, W18577, W15831, W15751);
nand G19248 (W17851, W15831, W18578);
nand G19249 (W17852, W15829, W18578);
nor G19250 (W17853, W18579, W18580);
not G19251 (W17854, W17856);
nor G19252 (W17855, W18581, W18582);
not G19253 (W17856, W18583);
nor G19254 (W17857, W18584, W18585);
not G19255 (W17858, W17860);
nor G19256 (W17859, W18586, W18587);
not G19257 (W17860, W18588);
not G19258 (W17861, W18589);
not G19259 (W17862, W18590);
not G19260 (W17863, W5385);
not G19261 (W17864, W18591);
not G19262 (W17865, W18592);
not G19263 (W17866, W18593);
not G19264 (W17867, W18594);
not G19265 (W17868, W18595);
and G19266 (W17869, W18596, W18597);
nand G19267 (W17870, I1365, I1366);
nand G19268 (W17871, I1367, I1368);
nand G19269 (W17872, I1369, I1370);
nand G19270 (W17873, I1371, I1372);
nand G19271 (W17874, I1373, I1374);
nand G19272 (W17875, I1375, I1376);
nand G19273 (W17876, I1377, I1378);
nand G19274 (W17877, I1379, I1380);
not G19275 (W17878, W18598);
and G19276 (W17879, W18599, W18600, W18601, W18602);
and G19277 (W17880, W18603, W18604, W18605);
and G19278 (W17881, W18606, W18607, W18608, W18609);
and G19279 (W17882, W18610, W18607, W18611, W18612);
and G19280 (W17883, W18607, W18611, W18613);
and G19281 (W17884, W18610, W18614, W18615);
and G19282 (W17885, W5253, W5252, W18606, W18614);
and G19283 (W17886, W18616, W5251, W18610, W18617);
and G19284 (W17887, W5250, W18610, W18607, W18608);
or G19285 (W17888, W18618, W18619, W18620);
and G19286 (W17889, W5253, W5251, W18617, W18608);
and G19287 (W17890, W5252, W18621, W18610, W18614);
and G19288 (W17891, W18616, W5251, W18622);
and G19289 (W17892, W5250, W18606, W18614);
and G19290 (W17893, W18617, W18608, W18623);
and G19291 (W17894, W18607, W18608, W18624);
or G19292 (W17895, W18625, W18626, W18627);
and G19293 (W17896, W18616, W18628, W18610, W18622);
and G19294 (W17897, W5253, W5250, W18606, W18611);
or G19295 (W17898, W18629, W18630, W18631);
and G19296 (W17899, W18632, W18633, W18634, W18635);
and G19297 (W17900, W18636, W18633, W18637, W18638);
and G19298 (W17901, W18633, W18637, W18639);
and G19299 (W17902, W18636, W18640, W18641);
and G19300 (W17903, W4978, W4977, W18632, W18640);
and G19301 (W17904, W18642, W4976, W18636, W18643);
and G19302 (W17905, W4975, W18636, W18633, W18634);
or G19303 (W17906, W18644, W18645, W18646);
and G19304 (W17907, W4978, W4976, W18643, W18634);
and G19305 (W17908, W4977, W18647, W18636, W18640);
and G19306 (W17909, W18642, W4976, W18648);
and G19307 (W17910, W4975, W18632, W18640);
and G19308 (W17911, W18643, W18634, W18649);
and G19309 (W17912, W18633, W18634, W18650);
or G19310 (W17913, W18651, W18652, W18653);
and G19311 (W17914, W18642, W18654, W18636, W18648);
and G19312 (W17915, W4978, W4975, W18632, W18637);
or G19313 (W17916, W18655, W18656, W18657);
and G19314 (W17917, W18658, W18659, W18660, W18661);
and G19315 (W17918, W18662, W18659, W18663, W18664);
and G19316 (W17919, W18659, W18663, W18665);
and G19317 (W17920, W18662, W18666, W18667);
and G19318 (W17921, W4703, W4702, W18658, W18666);
and G19319 (W17922, W18668, W4701, W18662, W18669);
and G19320 (W17923, W4700, W18662, W18659, W18660);
or G19321 (W17924, W18670, W18671, W18672);
and G19322 (W17925, W4703, W4701, W18669, W18660);
and G19323 (W17926, W4702, W18673, W18662, W18666);
and G19324 (W17927, W18668, W4701, W18674);
and G19325 (W17928, W4700, W18658, W18666);
and G19326 (W17929, W18669, W18660, W18675);
and G19327 (W17930, W18659, W18660, W18676);
or G19328 (W17931, W18677, W18678, W18679);
and G19329 (W17932, W18668, W18680, W18662, W18674);
and G19330 (W17933, W4703, W4700, W18658, W18663);
or G19331 (W17934, W18681, W18682, W18683);
and G19332 (W17935, W18684, W18685, W18686, W18687);
and G19333 (W17936, W18688, W18685, W18689, W18690);
and G19334 (W17937, W18685, W18689, W18691);
and G19335 (W17938, W18688, W18692, W18693);
and G19336 (W17939, W4428, W4427, W18684, W18692);
and G19337 (W17940, W18694, W4426, W18688, W18695);
and G19338 (W17941, W4425, W18688, W18685, W18686);
or G19339 (W17942, W18696, W18697, W18698);
and G19340 (W17943, W4428, W4426, W18695, W18686);
and G19341 (W17944, W4427, W18699, W18688, W18692);
and G19342 (W17945, W18694, W4426, W18700);
and G19343 (W17946, W4425, W18684, W18692);
and G19344 (W17947, W18695, W18686, W18701);
and G19345 (W17948, W18685, W18686, W18702);
or G19346 (W17949, W18703, W18704, W18705);
and G19347 (W17950, W18694, W18706, W18688, W18700);
and G19348 (W17951, W4428, W4425, W18684, W18689);
or G19349 (W17952, W18707, W18708, W18709);
not G19350 (W17953, W18710);
not G19351 (W17954, I1555);
not G19352 (W17955, I1531);
nand G19353 (W17956, W8442, W17957);
nand G19354 (W17957, W16588, W17983);
nand G19355 (W17958, W8432, W17959);
nand G19356 (W17959, W16588, W17981);
nor G19357 (W17960, W18711, W18712, W18713);
nand G19358 (W17961, W13835, W18714, W18715, W18716);
nand G19359 (W17962, W8432, W17963);
nand G19360 (W17963, W16588, W17985);
nand G19361 (W17964, W8442, W17965);
nand G19362 (W17965, W16588, W17327);
nand G19363 (W17966, W8432, W17967);
nand G19364 (W17967, W16588, W17991);
nand G19365 (W17968, W15125, W15113);
nand G19366 (W17969, W15133, W15129);
nand G19367 (W17970, W15107, W15098);
nand G19368 (W17971, W15094, W15103);
nand G19369 (W17972, W8442, W17973);
nand G19370 (W17973, W16588, W17989);
nand G19371 (W17974, W8432, W17975);
nand G19372 (W17975, W16588, W17325);
nand G19373 (W17976, W8442, W17977);
nand G19374 (W17977, W16588, W17993);
nor G19375 (W17978, W18717, W18718, W18719);
nor G19376 (W17979, W18720, W18721, W18722);
nand G19377 (W17980, W11992, W17981);
not G19378 (W17981, W18723);
nand G19379 (W17982, W11988, W17983);
not G19380 (W17983, W18724);
nand G19381 (W17984, W11986, W17985);
not G19382 (W17985, W18725);
nor G19383 (W17986, W18726, W18727, W18728);
nor G19384 (W17987, W18729, W18730, W18731);
nand G19385 (W17988, W12006, W17989);
not G19386 (W17989, W18732);
nand G19387 (W17990, W12004, W17991);
not G19388 (W17991, W18733);
nand G19389 (W17992, W12000, W17993);
not G19390 (W17993, W18734);
nand G19391 (W17994, W9009, W17995);
not G19392 (W17995, W18735);
nand G19393 (W17996, W9013, W17997);
not G19394 (W17997, W18736);
nand G19395 (W17998, W9033, W18737);
nand G19396 (W17999, W18738, W18737);
nand G19397 (W18000, W9041, W18739);
nand G19398 (W18001, W18740, W18739);
nand G19399 (W18002, W9005, W18741);
nand G19400 (W18003, W18742, W18741);
nand G19401 (W18004, W9029, W18005);
not G19402 (W18005, W18743);
nand G19403 (W18006, W9037, W18007);
not G19404 (W18007, W18744);
nand G19405 (W18008, W9017, W18745);
nand G19406 (W18009, W18746, W18745);
nand G19407 (W18010, W9021, W18747);
nand G19408 (W18011, W18748, W18747);
nand G19409 (W18012, W9025, W18749);
nand G19410 (W18013, W18750, W18749);
and G19411 (W18014, W13950, I650);
and G19412 (W18015, W13951, I651);
and G19413 (W18016, W9107, I652);
nand G19414 (W18017, W18751, W18752, W18753);
nor G19415 (W18018, W18754, W18755);
nor G19416 (W18019, W16057, W17356);
and G19417 (W18020, W17422, W13984);
and G19418 (W18021, W18756, W15243, W18757);
and G19419 (W18022, W15175, W12099, W18757);
and G19420 (W18023, W13950, I653);
and G19421 (W18024, W13951, I654);
and G19422 (W18025, W9107, I655);
nand G19423 (W18026, W18758, W18752, W18753, W18751);
not G19424 (W18027, W18759);
and G19425 (W18028, W13950, I656);
and G19426 (W18029, W13951, I657);
and G19427 (W18030, W9107, I658);
nand G19428 (W18031, W18047, W18760);
and G19429 (W18032, W13950, I659);
and G19430 (W18033, W13951, I660);
and G19431 (W18034, W9107, I661);
nor G19432 (W18035, W18055, W18761);
and G19433 (W18036, W13950, I663);
and G19434 (W18037, W13951, I664);
and G19435 (W18038, W9107, I662);
nor G19436 (W18039, W18059, W18762);
and G19437 (W18040, W13950, I667);
and G19438 (W18041, W13951, I665);
and G19439 (W18042, W9107, I666);
nor G19440 (W18043, W18017, W18763);
and G19441 (W18044, W13950, I668);
and G19442 (W18045, W13951, I669);
and G19443 (W18046, W9107, I670);
not G19444 (W18047, W18019);
and G19445 (W18048, W13950, I671);
and G19446 (W18049, W13951, I672);
and G19447 (W18050, W9107, I673);
nor G19448 (W18051, W18026, W18764);
and G19449 (W18052, W13950, I674);
and G19450 (W18053, W13951, I675);
and G19451 (W18054, W9107, I676);
not G19452 (W18055, W18752);
and G19453 (W18056, W13950, I677);
and G19454 (W18057, W13951, I678);
and G19455 (W18058, W9107, I679);
nand G19456 (W18059, W18753, W18752);
or G19457 (W18060, W15994, W13982);
or G19458 (W18061, W18765, W18766);
not G19459 (W18062, W12156);
nor G19460 (W18063, W18767, W18768);
not G19461 (W18064, W18065);
not G19462 (W18065, W18769);
and G19463 (W18066, W18770, W18771);
and G19464 (W18067, W18772, W18773);
not G19465 (W18068, W12156);
nand G19466 (W18069, W18774, W18775, W18776);
nand G19467 (W18070, W18777, W18778, W18779);
nand G19468 (W18071, W9108, W15194, W18780);
nand G19469 (W18072, I743, W16660);
nand G19470 (W18073, I744, W16688);
nand G19471 (W18074, I740, W18781);
nand G19472 (W18075, W16674, W18781);
nand G19473 (W18076, I741, W18782);
nand G19474 (W18077, W16652, W18782);
nand G19475 (W18078, I742, W18783);
nand G19476 (W18079, W16682, W18783);
nand G19477 (W18080, I748, W16645);
nand G19478 (W18081, I749, W16678);
nand G19479 (W18082, I745, W18784);
nand G19480 (W18083, W16666, W18784);
nand G19481 (W18084, I746, W18785);
nand G19482 (W18085, W16638, W18785);
nand G19483 (W18086, I747, W18786);
nand G19484 (W18087, W16670, W18786);
and G19485 (W18088, W13950, W9136);
and G19486 (W18089, W13951, W9133);
and G19487 (W18090, W9107, W9130);
not G19488 (W18091, W18787);
not G19489 (W18092, W18788);
not G19490 (W18093, W18789);
not G19491 (W18094, W18790);
not G19492 (W18095, W18791);
not G19493 (W18096, W18792);
not G19494 (W18097, W18793);
not G19495 (W18098, W18794);
not G19496 (W18099, W18795);
nand G19497 (W18100, W15263, W15261);
and G19498 (W18101, W18796, W18797);
not G19499 (W18102, W18798);
and G19500 (W18103, W18799, W18800);
and G19501 (W18104, W18801, W18802);
not G19502 (W18105, W15271);
and G19503 (W18106, W18803, W18804);
and G19504 (W18107, W18805, W18806);
and G19505 (W18108, W18807, W18808);
and G19506 (W18109, W18809, W18810);
not G19507 (W18110, W15271);
not G19508 (W18111, W18811);
nand G19509 (W18112, W18812, W16717);
not G19510 (W18113, I1556);
not G19511 (W18114, I1533);
nand G19512 (W18115, W9215, W18116);
nand G19513 (W18116, W16743, W18142);
nand G19514 (W18117, W9205, W18118);
nand G19515 (W18118, W16743, W18140);
nor G19516 (W18119, W18813, W18814, W18815);
nand G19517 (W18120, W14132, W18816, W18817, W18818);
nand G19518 (W18121, W9205, W18122);
nand G19519 (W18122, W16743, W18144);
nand G19520 (W18123, W9215, W18124);
nand G19521 (W18124, W16743, W17473);
nand G19522 (W18125, W9205, W18126);
nand G19523 (W18126, W16743, W18150);
nand G19524 (W18127, W15322, W15310);
nand G19525 (W18128, W15330, W15326);
nand G19526 (W18129, W15304, W15295);
nand G19527 (W18130, W15291, W15300);
nand G19528 (W18131, W9215, W18132);
nand G19529 (W18132, W16743, W18148);
nand G19530 (W18133, W9205, W18134);
nand G19531 (W18134, W16743, W17471);
nand G19532 (W18135, W9215, W18136);
nand G19533 (W18136, W16743, W18152);
nor G19534 (W18137, W18819, W18820, W18821);
nor G19535 (W18138, W18822, W18823, W18824);
nand G19536 (W18139, W12398, W18140);
not G19537 (W18140, W18825);
nand G19538 (W18141, W12394, W18142);
not G19539 (W18142, W18826);
nand G19540 (W18143, W12392, W18144);
not G19541 (W18144, W18827);
nor G19542 (W18145, W18828, W18829, W18830);
nor G19543 (W18146, W18831, W18832, W18833);
nand G19544 (W18147, W12412, W18148);
not G19545 (W18148, W18834);
nand G19546 (W18149, W12410, W18150);
not G19547 (W18150, W18835);
nand G19548 (W18151, W12406, W18152);
not G19549 (W18152, W18836);
nand G19550 (W18153, W9782, W18154);
not G19551 (W18154, W18837);
nand G19552 (W18155, W9786, W18156);
not G19553 (W18156, W18838);
nand G19554 (W18157, W9806, W18839);
nand G19555 (W18158, W18840, W18839);
nand G19556 (W18159, W9814, W18841);
nand G19557 (W18160, W18842, W18841);
nand G19558 (W18161, W9778, W18843);
nand G19559 (W18162, W18844, W18843);
nand G19560 (W18163, W9802, W18164);
not G19561 (W18164, W18845);
nand G19562 (W18165, W9810, W18166);
not G19563 (W18166, W18846);
nand G19564 (W18167, W9790, W18847);
nand G19565 (W18168, W18848, W18847);
nand G19566 (W18169, W9794, W18849);
nand G19567 (W18170, W18850, W18849);
nand G19568 (W18171, W9798, W18851);
nand G19569 (W18172, W18852, W18851);
and G19570 (W18173, W14244, I851);
and G19571 (W18174, W14245, I852);
and G19572 (W18175, W9880, I853);
nand G19573 (W18176, W18853, W18854, W18855);
nor G19574 (W18177, W18856, W18857);
nor G19575 (W18178, W16187, W17502);
and G19576 (W18179, W17568, W14278);
and G19577 (W18180, W18858, W15437, W18859);
and G19578 (W18181, W15369, W12505, W18859);
and G19579 (W18182, W14244, I854);
and G19580 (W18183, W14245, I855);
and G19581 (W18184, W9880, I856);
nand G19582 (W18185, W18860, W18854, W18855, W18853);
not G19583 (W18186, W18861);
and G19584 (W18187, W14244, I857);
and G19585 (W18188, W14245, I858);
and G19586 (W18189, W9880, I859);
nand G19587 (W18190, W18206, W18862);
and G19588 (W18191, W14244, I860);
and G19589 (W18192, W14245, I861);
and G19590 (W18193, W9880, I862);
nor G19591 (W18194, W18214, W18863);
and G19592 (W18195, W14244, I863);
and G19593 (W18196, W14245, I864);
and G19594 (W18197, W9880, I865);
nor G19595 (W18198, W18218, W18864);
and G19596 (W18199, W14244, I867);
and G19597 (W18200, W14245, I868);
and G19598 (W18201, W9880, I866);
nor G19599 (W18202, W18176, W18865);
and G19600 (W18203, W14244, I871);
and G19601 (W18204, W14245, I869);
and G19602 (W18205, W9880, I870);
not G19603 (W18206, W18178);
and G19604 (W18207, W14244, I874);
and G19605 (W18208, W14245, I872);
and G19606 (W18209, W9880, I873);
nor G19607 (W18210, W18185, W18866);
and G19608 (W18211, W14244, I875);
and G19609 (W18212, W14245, I876);
and G19610 (W18213, W9880, I877);
not G19611 (W18214, W18854);
and G19612 (W18215, W14244, I878);
and G19613 (W18216, W14245, I879);
and G19614 (W18217, W9880, I880);
nand G19615 (W18218, W18855, W18854);
or G19616 (W18219, W16124, W14276);
or G19617 (W18220, W18867, W18868);
not G19618 (W18221, W12562);
nor G19619 (W18222, W18869, W18870);
not G19620 (W18223, W18224);
not G19621 (W18224, W18871);
and G19622 (W18225, W18872, W18873);
and G19623 (W18226, W18874, W18875);
not G19624 (W18227, W12562);
nand G19625 (W18228, W18876, W18877, W18878);
nand G19626 (W18229, W18879, W18880, W18881);
nand G19627 (W18230, W9881, W15388, W18882);
nand G19628 (W18231, I944, W16815);
nand G19629 (W18232, I945, W16843);
nand G19630 (W18233, I941, W18883);
nand G19631 (W18234, W16829, W18883);
nand G19632 (W18235, I942, W18884);
nand G19633 (W18236, W16807, W18884);
nand G19634 (W18237, I943, W18885);
nand G19635 (W18238, W16837, W18885);
nand G19636 (W18239, I949, W16800);
nand G19637 (W18240, I950, W16833);
nand G19638 (W18241, I946, W18886);
nand G19639 (W18242, W16821, W18886);
nand G19640 (W18243, I947, W18887);
nand G19641 (W18244, W16793, W18887);
nand G19642 (W18245, I948, W18888);
nand G19643 (W18246, W16825, W18888);
and G19644 (W18247, W14244, W9909);
and G19645 (W18248, W14245, W9906);
and G19646 (W18249, W9880, W9903);
not G19647 (W18250, W18889);
not G19648 (W18251, W18890);
not G19649 (W18252, W18891);
not G19650 (W18253, W18892);
not G19651 (W18254, W18893);
not G19652 (W18255, W18894);
not G19653 (W18256, W18895);
not G19654 (W18257, W18896);
not G19655 (W18258, W18897);
nand G19656 (W18259, W15456, W15454);
and G19657 (W18260, W18898, W18899);
not G19658 (W18261, W18900);
and G19659 (W18262, W18901, W18902);
and G19660 (W18263, W18903, W18904);
not G19661 (W18264, W15464);
and G19662 (W18265, W18905, W18906);
and G19663 (W18266, W18907, W18908);
and G19664 (W18267, W18909, W18910);
and G19665 (W18268, W18911, W18912);
not G19666 (W18269, W15464);
not G19667 (W18270, W18913);
nand G19668 (W18271, W18914, W16872);
not G19669 (W18272, I1557);
not G19670 (W18273, I1535);
nand G19671 (W18274, W9988, W18275);
nand G19672 (W18275, W16898, W18301);
nand G19673 (W18276, W9978, W18277);
nand G19674 (W18277, W16898, W18299);
nor G19675 (W18278, W18915, W18916, W18917);
nand G19676 (W18279, W14425, W18918, W18919, W18920);
nand G19677 (W18280, W9978, W18281);
nand G19678 (W18281, W16898, W18303);
nand G19679 (W18282, W9988, W18283);
nand G19680 (W18283, W16898, W17619);
nand G19681 (W18284, W9978, W18285);
nand G19682 (W18285, W16898, W18309);
nand G19683 (W18286, W15515, W15503);
nand G19684 (W18287, W15523, W15519);
nand G19685 (W18288, W15497, W15488);
nand G19686 (W18289, W15484, W15493);
nand G19687 (W18290, W9988, W18291);
nand G19688 (W18291, W16898, W18307);
nand G19689 (W18292, W9978, W18293);
nand G19690 (W18293, W16898, W17617);
nand G19691 (W18294, W9988, W18295);
nand G19692 (W18295, W16898, W18311);
nor G19693 (W18296, W18921, W18922, W18923);
nor G19694 (W18297, W18924, W18925, W18926);
nand G19695 (W18298, W12804, W18299);
not G19696 (W18299, W18927);
nand G19697 (W18300, W12800, W18301);
not G19698 (W18301, W18928);
nand G19699 (W18302, W12798, W18303);
not G19700 (W18303, W18929);
nor G19701 (W18304, W18930, W18931, W18932);
nor G19702 (W18305, W18933, W18934, W18935);
nand G19703 (W18306, W12818, W18307);
not G19704 (W18307, W18936);
nand G19705 (W18308, W12816, W18309);
not G19706 (W18309, W18937);
nand G19707 (W18310, W12812, W18311);
not G19708 (W18311, W18938);
nand G19709 (W18312, W10551, W18313);
not G19710 (W18313, W18939);
nand G19711 (W18314, W10555, W18315);
not G19712 (W18315, W18940);
nand G19713 (W18316, W10575, W18941);
nand G19714 (W18317, W18942, W18941);
nand G19715 (W18318, W10583, W18943);
nand G19716 (W18319, W18944, W18943);
nand G19717 (W18320, W10587, W18945);
nand G19718 (W18321, W18946, W18945);
nand G19719 (W18322, W10571, W18323);
not G19720 (W18323, W18947);
nand G19721 (W18324, W10579, W18325);
not G19722 (W18325, W18948);
nand G19723 (W18326, W10559, W18949);
nand G19724 (W18327, W18950, W18949);
nand G19725 (W18328, W10563, W18951);
nand G19726 (W18329, W18952, W18951);
nand G19727 (W18330, W10567, W18953);
nand G19728 (W18331, W18954, W18953);
and G19729 (W18332, W14537, I1052);
and G19730 (W18333, W14538, I1053);
and G19731 (W18334, W10653, I1054);
nand G19732 (W18335, W18955, W18956, W18957);
nor G19733 (W18336, W18958, W18959);
nor G19734 (W18337, W16317, W17648);
and G19735 (W18338, W17714, W14571);
and G19736 (W18339, W18960, W15630, W18961);
and G19737 (W18340, W15562, W12911, W18961);
and G19738 (W18341, W14537, I1055);
and G19739 (W18342, W14538, I1056);
and G19740 (W18343, W10653, I1057);
nand G19741 (W18344, W18962, W18956, W18957, W18955);
not G19742 (W18345, W18963);
and G19743 (W18346, W14537, I1058);
and G19744 (W18347, W14538, I1059);
and G19745 (W18348, W10653, I1060);
nand G19746 (W18349, W18365, W18964);
and G19747 (W18350, W14537, I1061);
and G19748 (W18351, W14538, I1062);
and G19749 (W18352, W10653, I1063);
nor G19750 (W18353, W18373, W18965);
and G19751 (W18354, W14537, I1064);
and G19752 (W18355, W14538, I1065);
and G19753 (W18356, W10653, I1066);
nor G19754 (W18357, W18377, W18966);
and G19755 (W18358, W14537, I1067);
and G19756 (W18359, W14538, I1068);
and G19757 (W18360, W10653, I1069);
nor G19758 (W18361, W18335, W18967);
and G19759 (W18362, W14537, I1071);
and G19760 (W18363, W14538, I1072);
and G19761 (W18364, W10653, I1070);
not G19762 (W18365, W18337);
and G19763 (W18366, W14537, I1074);
and G19764 (W18367, W14538, I1075);
and G19765 (W18368, W10653, I1073);
nor G19766 (W18369, W18344, W18968);
and G19767 (W18370, W14537, I1078);
and G19768 (W18371, W14538, I1076);
and G19769 (W18372, W10653, I1077);
not G19770 (W18373, W18956);
and G19771 (W18374, W14537, I1079);
and G19772 (W18375, W14538, I1080);
and G19773 (W18376, W10653, I1081);
nand G19774 (W18377, W18957, W18956);
or G19775 (W18378, W16254, W14569);
or G19776 (W18379, W18969, W18970);
not G19777 (W18380, W12968);
nor G19778 (W18381, W18971, W18972);
not G19779 (W18382, W18383);
not G19780 (W18383, W18973);
and G19781 (W18384, W18974, W18975);
and G19782 (W18385, W18976, W18977);
not G19783 (W18386, W12968);
nand G19784 (W18387, W18978, W18979, W18980);
nand G19785 (W18388, W18981, W18982, W18983);
nand G19786 (W18389, W10654, W15581, W18984);
nand G19787 (W18390, I1145, W16970);
nand G19788 (W18391, I1146, W16998);
nand G19789 (W18392, I1142, W18985);
nand G19790 (W18393, W16984, W18985);
nand G19791 (W18394, I1143, W18986);
nand G19792 (W18395, W16962, W18986);
nand G19793 (W18396, I1144, W18987);
nand G19794 (W18397, W16992, W18987);
nand G19795 (W18398, I1150, W16955);
nand G19796 (W18399, I1151, W16988);
nand G19797 (W18400, I1147, W18988);
nand G19798 (W18401, W16976, W18988);
nand G19799 (W18402, I1148, W18989);
nand G19800 (W18403, W16948, W18989);
nand G19801 (W18404, I1149, W18990);
nand G19802 (W18405, W16980, W18990);
and G19803 (W18406, W14537, W10682);
and G19804 (W18407, W14538, W10679);
and G19805 (W18408, W10653, W10676);
not G19806 (W18409, W18991);
not G19807 (W18410, W18992);
not G19808 (W18411, W18993);
not G19809 (W18412, W18994);
not G19810 (W18413, W18995);
not G19811 (W18414, W18996);
not G19812 (W18415, W18997);
not G19813 (W18416, W18998);
not G19814 (W18417, W18999);
nand G19815 (W18418, W15649, W15647);
and G19816 (W18419, W19000, W19001);
not G19817 (W18420, W19002);
and G19818 (W18421, W19003, W19004);
and G19819 (W18422, W19005, W19006);
not G19820 (W18423, W15657);
and G19821 (W18424, W19007, W19008);
and G19822 (W18425, W19009, W19010);
and G19823 (W18426, W19011, W19012);
and G19824 (W18427, W19013, W19014);
not G19825 (W18428, W15657);
not G19826 (W18429, W19015);
nand G19827 (W18430, W19016, W17027);
not G19828 (W18431, I1558);
not G19829 (W18432, W11015);
not G19830 (W18433, I1537);
nand G19831 (W18434, W10761, W18435);
nand G19832 (W18435, W17053, W18461);
nand G19833 (W18436, W10751, W18437);
nand G19834 (W18437, W17053, W18459);
nor G19835 (W18438, W19017, W19018, W19019);
nand G19836 (W18439, W14718, W19020, W19021, W19022);
nand G19837 (W18440, W10751, W18441);
nand G19838 (W18441, W17053, W18463);
nand G19839 (W18442, W10761, W18443);
nand G19840 (W18443, W17053, W17766);
nand G19841 (W18444, W10751, W18445);
nand G19842 (W18445, W17053, W18469);
nand G19843 (W18446, W15708, W15696);
nand G19844 (W18447, W15716, W15712);
nand G19845 (W18448, W15690, W15681);
nand G19846 (W18449, W15677, W15686);
nand G19847 (W18450, W10761, W18451);
nand G19848 (W18451, W17053, W18467);
nand G19849 (W18452, W10751, W18453);
nand G19850 (W18453, W17053, W17764);
nand G19851 (W18454, W10761, W18455);
nand G19852 (W18455, W17053, W18471);
nor G19853 (W18456, W19023, W19024, W19025);
nor G19854 (W18457, W19026, W19027, W19028);
nand G19855 (W18458, W13210, W18459);
not G19856 (W18459, W19029);
nand G19857 (W18460, W13206, W18461);
not G19858 (W18461, W19030);
nand G19859 (W18462, W13204, W18463);
not G19860 (W18463, W19031);
nor G19861 (W18464, W19032, W19033, W19034);
nor G19862 (W18465, W19035, W19036, W19037);
nand G19863 (W18466, W13224, W18467);
not G19864 (W18467, W19038);
nand G19865 (W18468, W13222, W18469);
not G19866 (W18469, W19039);
nand G19867 (W18470, W13218, W18471);
not G19868 (W18471, W19040);
nand G19869 (W18472, W11363, W18473);
not G19870 (W18473, W19041);
nand G19871 (W18474, W11324, W18475);
not G19872 (W18475, W19042);
nand G19873 (W18476, W11344, W19043);
nand G19874 (W18477, W19044, W19043);
nand G19875 (W18478, W11352, W19045);
nand G19876 (W18479, W19046, W19045);
nand G19877 (W18480, W11356, W19047);
nand G19878 (W18481, W19048, W19047);
nand G19879 (W18482, W11340, W18483);
not G19880 (W18483, W19049);
nand G19881 (W18484, W11348, W18485);
not G19882 (W18485, W19050);
nand G19883 (W18486, W11328, W19051);
nand G19884 (W18487, W19052, W19051);
nand G19885 (W18488, W11332, W19053);
nand G19886 (W18489, W19054, W19053);
nand G19887 (W18490, W11336, W19055);
nand G19888 (W18491, W19056, W19055);
and G19889 (W18492, W14808, I1253);
and G19890 (W18493, W14809, I1254);
and G19891 (W18494, W11426, I1255);
nand G19892 (W18495, W19057, W19058, W19059);
nor G19893 (W18496, W19060, W19061);
nor G19894 (W18497, W16459, W17795);
and G19895 (W18498, W17861, W14842);
and G19896 (W18499, W19062, W15812, W19063);
and G19897 (W18500, W15750, W13306, W19063);
and G19898 (W18501, W14808, I1256);
and G19899 (W18502, W14809, I1257);
and G19900 (W18503, W11426, I1258);
nand G19901 (W18504, W19064, W19058, W19059, W19057);
not G19902 (W18505, W19065);
and G19903 (W18506, W14808, I1259);
and G19904 (W18507, W14809, I1260);
and G19905 (W18508, W11426, I1261);
nand G19906 (W18509, W18525, W19066);
and G19907 (W18510, W14808, I1262);
and G19908 (W18511, W14809, I1263);
and G19909 (W18512, W11426, I1264);
nor G19910 (W18513, W18533, W19067);
and G19911 (W18514, W14808, I1265);
and G19912 (W18515, W14809, I1266);
and G19913 (W18516, W11426, I1267);
nor G19914 (W18517, W18537, W19068);
and G19915 (W18518, W14808, I1268);
and G19916 (W18519, W14809, I1269);
and G19917 (W18520, W11426, I1270);
nor G19918 (W18521, W18495, W19069);
and G19919 (W18522, W14808, I1271);
and G19920 (W18523, W14809, I1272);
and G19921 (W18524, W11426, I1273);
not G19922 (W18525, W18497);
and G19923 (W18526, W14808, I1274);
and G19924 (W18527, W14809, I1275);
and G19925 (W18528, W11426, I1276);
nor G19926 (W18529, W18504, W19070);
and G19927 (W18530, W14808, I1278);
and G19928 (W18531, W14809, I1279);
and G19929 (W18532, W11426, I1277);
not G19930 (W18533, W19058);
and G19931 (W18534, W14808, I1282);
and G19932 (W18535, W14809, I1280);
and G19933 (W18536, W11426, I1281);
nand G19934 (W18537, W19059, W19058);
or G19935 (W18538, W16390, W14840);
or G19936 (W18539, W19071, W19072);
not G19937 (W18540, W13363);
nor G19938 (W18541, W19073, W19074);
not G19939 (W18542, W18543);
not G19940 (W18543, W19075);
and G19941 (W18544, W19076, W19077);
and G19942 (W18545, W19078, W19079);
not G19943 (W18546, W13363);
nand G19944 (W18547, W19080, W19081, W19082);
nand G19945 (W18548, W19083, W19084, W19085);
nand G19946 (W18549, W11427, W15763, W19086);
nand G19947 (W18550, I1346, W17125);
nand G19948 (W18551, I1347, W17153);
nand G19949 (W18552, I1343, W19087);
nand G19950 (W18553, W17139, W19087);
nand G19951 (W18554, I1344, W19088);
nand G19952 (W18555, W17117, W19088);
nand G19953 (W18556, I1345, W19089);
nand G19954 (W18557, W17147, W19089);
nand G19955 (W18558, I1351, W17110);
nand G19956 (W18559, I1352, W17143);
nand G19957 (W18560, I1348, W19090);
nand G19958 (W18561, W17131, W19090);
nand G19959 (W18562, I1349, W19091);
nand G19960 (W18563, W17103, W19091);
nand G19961 (W18564, I1350, W19092);
nand G19962 (W18565, W17135, W19092);
and G19963 (W18566, W14808, W11455);
and G19964 (W18567, W14809, W11452);
and G19965 (W18568, W11426, W11449);
not G19966 (W18569, W19093);
not G19967 (W18570, W19094);
not G19968 (W18571, W19095);
not G19969 (W18572, W19096);
not G19970 (W18573, W19097);
not G19971 (W18574, W19098);
not G19972 (W18575, W19099);
not G19973 (W18576, W19100);
not G19974 (W18577, W19101);
nand G19975 (W18578, W15831, W15829);
and G19976 (W18579, W19102, W19103);
not G19977 (W18580, W19104);
and G19978 (W18581, W19105, W19106);
and G19979 (W18582, W19107, W19108);
not G19980 (W18583, W15839);
and G19981 (W18584, W19109, W19110);
and G19982 (W18585, W19111, W19112);
and G19983 (W18586, W19113, W19114);
and G19984 (W18587, W19115, W19116);
not G19985 (W18588, W15839);
not G19986 (W18589, W19117);
nand G19987 (W18590, W19118, W17182);
and G19988 (W18591, W19119, W19120, W19121, W19122);
and G19989 (W18592, W19123, W19124, W19125, W19126);
nor G19990 (W18593, W19127, W19128);
nor G19991 (W18594, W19129, W19130);
nor G19992 (W18595, W19131, W19132);
not G19993 (W18596, I1559);
not G19994 (W18597, W19133);
not G19995 (W18598, W19134);
nor G19996 (W18599, W19135, W19136, W19137);
nor G19997 (W18600, W19138, W19139, W19140);
nor G19998 (W18601, W19141, W19142, W19143);
and G19999 (W18602, W19144, W19145, W19146);
nor G20000 (W18603, W19147, W19148);
nor G20001 (W18604, W19149, W19150, W19151);
nor G20002 (W18605, W19152, W19153, W19154);
not G20003 (W18606, W19155);
not G20004 (W18607, W19156);
not G20005 (W18608, W19157);
and G20006 (W18609, W5253, W19158, W18628);
not G20007 (W18610, W19159);
not G20008 (W18611, W19160);
and G20009 (W18612, W18616, W19158, W18621);
and G20010 (W18613, W5253, W5251, W18606);
not G20011 (W18614, W19161);
and G20012 (W18615, W18616, W19158, W18628);
not G20013 (W18616, W5253);
not G20014 (W18617, W19162);
and G20015 (W18618, W5253, W19158, W18621, W18622);
and G20016 (W18619, W18616, W5252, W18617, W18608);
and G20017 (W18620, W5252, W18621, W18606, W18617);
not G20018 (W18621, W5251);
not G20019 (W18622, W19163);
and G20020 (W18623, W5253, W18628, W18610);
and G20021 (W18624, W18616, W5251, W18610);
and G20022 (W18625, W18607, W18608, W19164);
and G20023 (W18626, W18607, W18611, W19165);
and G20024 (W18627, W5253, W19158, W18606, W18617);
not G20025 (W18628, W5250);
and G20026 (W18629, W18607, W18614, W19166);
and G20027 (W18630, W5252, W18610, W18607, W18614);
and G20028 (W18631, W5253, W5251, W18610, W18617);
not G20029 (W18632, W19167);
not G20030 (W18633, W19168);
not G20031 (W18634, W19169);
and G20032 (W18635, W4978, W19170, W18654);
not G20033 (W18636, W19171);
not G20034 (W18637, W19172);
and G20035 (W18638, W18642, W19170, W18647);
and G20036 (W18639, W4978, W4976, W18632);
not G20037 (W18640, W19173);
and G20038 (W18641, W18642, W19170, W18654);
not G20039 (W18642, W4978);
not G20040 (W18643, W19174);
and G20041 (W18644, W4978, W19170, W18647, W18648);
and G20042 (W18645, W18642, W4977, W18643, W18634);
and G20043 (W18646, W4977, W18647, W18632, W18643);
not G20044 (W18647, W4976);
not G20045 (W18648, W19175);
and G20046 (W18649, W4978, W18654, W18636);
and G20047 (W18650, W18642, W4976, W18636);
and G20048 (W18651, W18633, W18634, W19176);
and G20049 (W18652, W18633, W18637, W19177);
and G20050 (W18653, W4978, W19170, W18632, W18643);
not G20051 (W18654, W4975);
and G20052 (W18655, W18633, W18640, W19178);
and G20053 (W18656, W4977, W18636, W18633, W18640);
and G20054 (W18657, W4978, W4976, W18636, W18643);
not G20055 (W18658, W19179);
not G20056 (W18659, W19180);
not G20057 (W18660, W19181);
and G20058 (W18661, W4703, W19182, W18680);
not G20059 (W18662, W19183);
not G20060 (W18663, W19184);
and G20061 (W18664, W18668, W19182, W18673);
and G20062 (W18665, W4703, W4701, W18658);
not G20063 (W18666, W19185);
and G20064 (W18667, W18668, W19182, W18680);
not G20065 (W18668, W4703);
not G20066 (W18669, W19186);
and G20067 (W18670, W4703, W19182, W18673, W18674);
and G20068 (W18671, W18668, W4702, W18669, W18660);
and G20069 (W18672, W4702, W18673, W18658, W18669);
not G20070 (W18673, W4701);
not G20071 (W18674, W19187);
and G20072 (W18675, W4703, W18680, W18662);
and G20073 (W18676, W18668, W4701, W18662);
and G20074 (W18677, W18659, W18660, W19188);
and G20075 (W18678, W18659, W18663, W19189);
and G20076 (W18679, W4703, W19182, W18658, W18669);
not G20077 (W18680, W4700);
and G20078 (W18681, W18659, W18666, W19190);
and G20079 (W18682, W4702, W18662, W18659, W18666);
and G20080 (W18683, W4703, W4701, W18662, W18669);
not G20081 (W18684, W19191);
not G20082 (W18685, W19192);
not G20083 (W18686, W19193);
and G20084 (W18687, W4428, W19194, W18706);
not G20085 (W18688, W19195);
not G20086 (W18689, W19196);
and G20087 (W18690, W18694, W19194, W18699);
and G20088 (W18691, W4428, W4426, W18684);
not G20089 (W18692, W19197);
and G20090 (W18693, W18694, W19194, W18706);
not G20091 (W18694, W4428);
not G20092 (W18695, W19198);
and G20093 (W18696, W4428, W19194, W18699, W18700);
and G20094 (W18697, W18694, W4427, W18695, W18686);
and G20095 (W18698, W4427, W18699, W18684, W18695);
not G20096 (W18699, W4426);
not G20097 (W18700, W19199);
and G20098 (W18701, W4428, W18706, W18688);
and G20099 (W18702, W18694, W4426, W18688);
and G20100 (W18703, W18685, W18686, W19200);
and G20101 (W18704, W18685, W18689, W19201);
and G20102 (W18705, W4428, W19194, W18684, W18695);
not G20103 (W18706, W4425);
and G20104 (W18707, W18685, W18692, W19202);
and G20105 (W18708, W4427, W18688, W18685, W18692);
and G20106 (W18709, W4428, W4426, W18688, W18695);
not G20107 (W18710, I1560);
and G20108 (W18711, W15138, W8430);
and G20109 (W18712, W8544, W8427);
and G20110 (W18713, W13643, W8424);
not G20111 (W18714, W19203);
and G20112 (W18715, W17325, W19204, W19205);
and G20113 (W18716, W17315, W17317, W19206);
and G20114 (W18717, W15138, W8468);
and G20115 (W18718, W8544, W8465);
and G20116 (W18719, W13643, W8462);
and G20117 (W18720, W15138, W8459);
and G20118 (W18721, W8544, W8456);
and G20119 (W18722, W13643, W8453);
nor G20120 (W18723, W19207, W19208, W19209);
nor G20121 (W18724, W19210, W19211, W19212);
nor G20122 (W18725, W19213, W19214, W19215);
and G20123 (W18726, W15138, W8513);
and G20124 (W18727, W8544, W8510);
and G20125 (W18728, W13643, W8507);
and G20126 (W18729, W15138, W8504);
and G20127 (W18730, W8544, W8501);
and G20128 (W18731, W13643, W8498);
nor G20129 (W18732, W19216, W19217, W19218);
nor G20130 (W18733, W19219, W19220, W19221);
nor G20131 (W18734, W19222, W19223, W19224);
nor G20132 (W18735, W19225, W19226, W19227);
nor G20133 (W18736, W19228, W19229, W19230);
nand G20134 (W18737, W9033, W18738);
not G20135 (W18738, W19231);
nand G20136 (W18739, W9041, W18740);
not G20137 (W18740, W19232);
nand G20138 (W18741, W9005, W18742);
not G20139 (W18742, W19233);
nor G20140 (W18743, W19234, W19235, W19236);
nor G20141 (W18744, W19237, W19238, W19239);
nand G20142 (W18745, W9017, W18746);
not G20143 (W18746, W19240);
nand G20144 (W18747, W9021, W18748);
not G20145 (W18748, W19241);
nand G20146 (W18749, W9025, W18750);
not G20147 (W18750, W19242);
nor G20148 (W18751, W18762, W19243);
nor G20149 (W18752, W18031, W19244);
nor G20150 (W18753, W18761, W19245);
and G20151 (W18754, W16058, W19246);
and G20152 (W18755, W19247, W19248);
nor G20153 (W18756, W15244, W15994, W12156);
not G20154 (W18757, W19249);
nor G20155 (W18758, W18763, W19250);
nor G20156 (W18759, W15244, W13983, W13984);
nor G20157 (W18760, W19251, W19252);
nor G20158 (W18761, W19253, W19254);
nor G20159 (W18762, W19255, W19256);
nor G20160 (W18763, W19257, W19258);
nor G20161 (W18764, W19259, W19260);
not G20162 (W18765, W17389);
not G20163 (W18766, W17388);
and G20164 (W18767, W19261, W19262);
and G20165 (W18768, W19263, W19264);
not G20166 (W18769, W12156);
nor G20167 (W18770, W19265, W19266);
not G20168 (W18771, W18773);
nor G20169 (W18772, W19267, W19268);
not G20170 (W18773, W19269);
nand G20171 (W18774, W19270, W19271, W19272);
nand G20172 (W18775, W19273, W19274, W19275);
nand G20173 (W18776, W19276, W19277, W19278);
nand G20174 (W18777, W19279, W19280, W19281);
nand G20175 (W18778, W19282, W19283, W19284);
nand G20176 (W18779, W19285, W19286, W19287);
not G20177 (W18780, W19288);
nand G20178 (W18781, I740, W16674);
nand G20179 (W18782, I741, W16652);
nand G20180 (W18783, I742, W16682);
nand G20181 (W18784, I745, W16666);
nand G20182 (W18785, I746, W16638);
nand G20183 (W18786, I747, W16670);
not G20184 (W18787, I223);
not G20185 (W18788, I224);
not G20186 (W18789, I225);
not G20187 (W18790, I226);
not G20188 (W18791, I227);
not G20189 (W18792, I228);
not G20190 (W18793, I229);
not G20191 (W18794, I230);
not G20192 (W18795, W16064);
nand G20193 (W18796, W17422, W18805);
not G20194 (W18797, W19289);
not G20195 (W18798, W19289);
nand G20196 (W18799, W18805, W19290);
not G20197 (W18800, W18802);
nand G20198 (W18801, W15274, W16732);
not G20199 (W18802, W19291);
nand G20200 (W18803, W18111, W18805);
not G20201 (W18804, W18806);
not G20202 (W18805, W18112);
not G20203 (W18806, W19292);
nor G20204 (W18807, W15274, W17422, W16732);
not G20205 (W18808, W18810);
nor G20206 (W18809, W15274, W18805);
not G20207 (W18810, W19293);
nor G20208 (W18811, W12257, W15194);
and G20209 (W18812, W9037, W9029);
and G20210 (W18813, W15335, W9203);
and G20211 (W18814, W9317, W9200);
and G20212 (W18815, W13642, W9197);
not G20213 (W18816, W19294);
and G20214 (W18817, W17471, W19295, W19296);
and G20215 (W18818, W17461, W17463, W19297);
and G20216 (W18819, W15335, W9241);
and G20217 (W18820, W9317, W9238);
and G20218 (W18821, W13642, W9235);
and G20219 (W18822, W15335, W9232);
and G20220 (W18823, W9317, W9229);
and G20221 (W18824, W13642, W9226);
nor G20222 (W18825, W19298, W19299, W19300);
nor G20223 (W18826, W19301, W19302, W19303);
nor G20224 (W18827, W19304, W19305, W19306);
and G20225 (W18828, W15335, W9286);
and G20226 (W18829, W9317, W9283);
and G20227 (W18830, W13642, W9280);
and G20228 (W18831, W15335, W9277);
and G20229 (W18832, W9317, W9274);
and G20230 (W18833, W13642, W9271);
nor G20231 (W18834, W19307, W19308, W19309);
nor G20232 (W18835, W19310, W19311, W19312);
nor G20233 (W18836, W19313, W19314, W19315);
nor G20234 (W18837, W19316, W19317, W19318);
nor G20235 (W18838, W19319, W19320, W19321);
nand G20236 (W18839, W9806, W18840);
not G20237 (W18840, W19322);
nand G20238 (W18841, W9814, W18842);
not G20239 (W18842, W19323);
nand G20240 (W18843, W9778, W18844);
not G20241 (W18844, W19324);
nor G20242 (W18845, W19325, W19326, W19327);
nor G20243 (W18846, W19328, W19329, W19330);
nand G20244 (W18847, W9790, W18848);
not G20245 (W18848, W19331);
nand G20246 (W18849, W9794, W18850);
not G20247 (W18850, W19332);
nand G20248 (W18851, W9798, W18852);
not G20249 (W18852, W19333);
nor G20250 (W18853, W18864, W19334);
nor G20251 (W18854, W18190, W19335);
nor G20252 (W18855, W18863, W19336);
and G20253 (W18856, W16188, W19337);
and G20254 (W18857, W19338, W19339);
nor G20255 (W18858, W15438, W16124, W12562);
not G20256 (W18859, W19340);
nor G20257 (W18860, W18865, W19341);
nor G20258 (W18861, W15438, W14277, W14278);
nor G20259 (W18862, W19342, W19343);
nor G20260 (W18863, W19344, W19345);
nor G20261 (W18864, W19346, W19347);
nor G20262 (W18865, W19348, W19349);
nor G20263 (W18866, W19350, W19351);
not G20264 (W18867, W17535);
not G20265 (W18868, W17534);
and G20266 (W18869, W19352, W19353);
and G20267 (W18870, W19354, W19355);
not G20268 (W18871, W12562);
nor G20269 (W18872, W19356, W19357);
not G20270 (W18873, W18875);
nor G20271 (W18874, W19358, W19359);
not G20272 (W18875, W19360);
nand G20273 (W18876, W19361, W19362, W19363);
nand G20274 (W18877, W19364, W19365, W19366);
nand G20275 (W18878, W19367, W19368, W19369);
nand G20276 (W18879, W19370, W19371, W19372);
nand G20277 (W18880, W19373, W19374, W19375);
nand G20278 (W18881, W19376, W19377, W19378);
not G20279 (W18882, W19379);
nand G20280 (W18883, I941, W16829);
nand G20281 (W18884, I942, W16807);
nand G20282 (W18885, I943, W16837);
nand G20283 (W18886, I946, W16821);
nand G20284 (W18887, I947, W16793);
nand G20285 (W18888, I948, W16825);
not G20286 (W18889, I247);
not G20287 (W18890, I248);
not G20288 (W18891, I249);
not G20289 (W18892, I250);
not G20290 (W18893, I251);
not G20291 (W18894, I252);
not G20292 (W18895, I253);
not G20293 (W18896, I254);
not G20294 (W18897, W16194);
nand G20295 (W18898, W17568, W18907);
not G20296 (W18899, W19380);
not G20297 (W18900, W19380);
nand G20298 (W18901, W18907, W19381);
not G20299 (W18902, W18904);
nand G20300 (W18903, W15467, W16887);
not G20301 (W18904, W19382);
nand G20302 (W18905, W18270, W18907);
not G20303 (W18906, W18908);
not G20304 (W18907, W18271);
not G20305 (W18908, W19383);
nor G20306 (W18909, W15467, W17568, W16887);
not G20307 (W18910, W18912);
nor G20308 (W18911, W15467, W18907);
not G20309 (W18912, W19384);
nor G20310 (W18913, W12663, W15388);
and G20311 (W18914, W9810, W9802);
and G20312 (W18915, W15528, W9976);
and G20313 (W18916, W10090, W9973);
and G20314 (W18917, W13641, W9970);
not G20315 (W18918, W19385);
and G20316 (W18919, W17617, W19386, W19387);
and G20317 (W18920, W17607, W17609, W19388);
and G20318 (W18921, W15528, W10014);
and G20319 (W18922, W10090, W10011);
and G20320 (W18923, W13641, W10008);
and G20321 (W18924, W15528, W10005);
and G20322 (W18925, W10090, W10002);
and G20323 (W18926, W13641, W9999);
nor G20324 (W18927, W19389, W19390, W19391);
nor G20325 (W18928, W19392, W19393, W19394);
nor G20326 (W18929, W19395, W19396, W19397);
and G20327 (W18930, W15528, W10059);
and G20328 (W18931, W10090, W10056);
and G20329 (W18932, W13641, W10053);
and G20330 (W18933, W15528, W10050);
and G20331 (W18934, W10090, W10047);
and G20332 (W18935, W13641, W10044);
nor G20333 (W18936, W19398, W19399, W19400);
nor G20334 (W18937, W19401, W19402, W19403);
nor G20335 (W18938, W19404, W19405, W19406);
nor G20336 (W18939, W19407, W19408, W19409);
nor G20337 (W18940, W19410, W19411, W19412);
nand G20338 (W18941, W10575, W18942);
not G20339 (W18942, W19413);
nand G20340 (W18943, W10583, W18944);
not G20341 (W18944, W19414);
nand G20342 (W18945, W10587, W18946);
not G20343 (W18946, W19415);
nor G20344 (W18947, W19416, W19417, W19418);
nor G20345 (W18948, W19419, W19420, W19421);
nand G20346 (W18949, W10559, W18950);
not G20347 (W18950, W19422);
nand G20348 (W18951, W10563, W18952);
not G20349 (W18952, W19423);
nand G20350 (W18953, W10567, W18954);
not G20351 (W18954, W19424);
nor G20352 (W18955, W18966, W19425);
nor G20353 (W18956, W18349, W19426);
nor G20354 (W18957, W18965, W19427);
and G20355 (W18958, W16318, W19428);
and G20356 (W18959, W19429, W19430);
nor G20357 (W18960, W15631, W16254, W12968);
not G20358 (W18961, W19431);
nor G20359 (W18962, W18967, W19432);
nor G20360 (W18963, W15631, W14570, W14571);
nor G20361 (W18964, W19433, W19434);
nor G20362 (W18965, W19435, W19436);
nor G20363 (W18966, W19437, W19438);
nor G20364 (W18967, W19439, W19440);
nor G20365 (W18968, W19441, W19442);
not G20366 (W18969, W17681);
not G20367 (W18970, W17680);
and G20368 (W18971, W19443, W19444);
and G20369 (W18972, W19445, W19446);
not G20370 (W18973, W12968);
nor G20371 (W18974, W19447, W19448);
not G20372 (W18975, W18977);
nor G20373 (W18976, W19449, W19450);
not G20374 (W18977, W19451);
nand G20375 (W18978, W19452, W19453, W19454);
nand G20376 (W18979, W19455, W19456, W19457);
nand G20377 (W18980, W19458, W19459, W19460);
nand G20378 (W18981, W19461, W19462, W19463);
nand G20379 (W18982, W19464, W19465, W19466);
nand G20380 (W18983, W19467, W19468, W19469);
not G20381 (W18984, W19470);
nand G20382 (W18985, I1142, W16984);
nand G20383 (W18986, I1143, W16962);
nand G20384 (W18987, I1144, W16992);
nand G20385 (W18988, I1147, W16976);
nand G20386 (W18989, I1148, W16948);
nand G20387 (W18990, I1149, W16980);
not G20388 (W18991, I239);
not G20389 (W18992, I240);
not G20390 (W18993, I241);
not G20391 (W18994, I242);
not G20392 (W18995, I243);
not G20393 (W18996, I244);
not G20394 (W18997, I245);
not G20395 (W18998, I246);
not G20396 (W18999, W16324);
nand G20397 (W19000, W17714, W19009);
not G20398 (W19001, W19471);
not G20399 (W19002, W19471);
nand G20400 (W19003, W19009, W19472);
not G20401 (W19004, W19006);
nand G20402 (W19005, W15660, W17042);
not G20403 (W19006, W19473);
nand G20404 (W19007, W18429, W19009);
not G20405 (W19008, W19010);
not G20406 (W19009, W18430);
not G20407 (W19010, W19474);
nor G20408 (W19011, W15660, W17714, W17042);
not G20409 (W19012, W19014);
nor G20410 (W19013, W15660, W19009);
not G20411 (W19014, W19475);
nor G20412 (W19015, W13069, W15581);
and G20413 (W19016, W10579, W10571);
and G20414 (W19017, W15721, W10749);
and G20415 (W19018, W10863, W10746);
and G20416 (W19019, W13640, W10743);
not G20417 (W19020, W19476);
and G20418 (W19021, W17764, W19477, W19478);
and G20419 (W19022, W17754, W17756, W19479);
and G20420 (W19023, W15721, W10787);
and G20421 (W19024, W10863, W10784);
and G20422 (W19025, W13640, W10781);
and G20423 (W19026, W15721, W10778);
and G20424 (W19027, W10863, W10775);
and G20425 (W19028, W13640, W10772);
nor G20426 (W19029, W19480, W19481, W19482);
nor G20427 (W19030, W19483, W19484, W19485);
nor G20428 (W19031, W19486, W19487, W19488);
and G20429 (W19032, W15721, W10832);
and G20430 (W19033, W10863, W10829);
and G20431 (W19034, W13640, W10826);
and G20432 (W19035, W15721, W10823);
and G20433 (W19036, W10863, W10820);
and G20434 (W19037, W13640, W10817);
nor G20435 (W19038, W19489, W19490, W19491);
nor G20436 (W19039, W19492, W19493, W19494);
nor G20437 (W19040, W19495, W19496, W19497);
nor G20438 (W19041, W19498, W19499, W19500);
nor G20439 (W19042, W19501, W19502, W19503);
nand G20440 (W19043, W11344, W19044);
not G20441 (W19044, W19504);
nand G20442 (W19045, W11352, W19046);
not G20443 (W19046, W19505);
nand G20444 (W19047, W11356, W19048);
not G20445 (W19048, W19506);
nor G20446 (W19049, W19507, W19508, W19509);
nor G20447 (W19050, W19510, W19511, W19512);
nand G20448 (W19051, W11328, W19052);
not G20449 (W19052, W19513);
nand G20450 (W19053, W11332, W19054);
not G20451 (W19054, W19514);
nand G20452 (W19055, W11336, W19056);
not G20453 (W19056, W19515);
nor G20454 (W19057, W19068, W19516);
nor G20455 (W19058, W18509, W19517);
nor G20456 (W19059, W19067, W19518);
and G20457 (W19060, W16460, W19519);
and G20458 (W19061, W19520, W19521);
nor G20459 (W19062, W15813, W16390, W13363);
not G20460 (W19063, W19522);
nor G20461 (W19064, W19069, W19523);
nor G20462 (W19065, W15813, W14841, W14842);
nor G20463 (W19066, W19524, W19525);
nor G20464 (W19067, W19526, W19527);
nor G20465 (W19068, W19528, W19529);
nor G20466 (W19069, W19530, W19531);
nor G20467 (W19070, W19532, W19533);
not G20468 (W19071, W17828);
not G20469 (W19072, W17827);
and G20470 (W19073, W19534, W19535);
and G20471 (W19074, W19536, W19537);
not G20472 (W19075, W13363);
nor G20473 (W19076, W19538, W19539);
not G20474 (W19077, W19079);
nor G20475 (W19078, W19540, W19541);
not G20476 (W19079, W19542);
nand G20477 (W19080, W19543, W19544, W19545);
nand G20478 (W19081, W19546, W19547, W19548);
nand G20479 (W19082, W19549, W19550, W19551);
nand G20480 (W19083, W19552, W19553, W19554);
nand G20481 (W19084, W19555, W19556, W19557);
nand G20482 (W19085, W19558, W19559, W19560);
not G20483 (W19086, W19561);
nand G20484 (W19087, I1343, W17139);
nand G20485 (W19088, I1344, W17117);
nand G20486 (W19089, I1345, W17147);
nand G20487 (W19090, I1348, W17131);
nand G20488 (W19091, I1349, W17103);
nand G20489 (W19092, I1350, W17135);
not G20490 (W19093, I231);
not G20491 (W19094, I232);
not G20492 (W19095, I233);
not G20493 (W19096, I234);
not G20494 (W19097, I235);
not G20495 (W19098, I236);
not G20496 (W19099, I237);
not G20497 (W19100, I238);
not G20498 (W19101, W16466);
nand G20499 (W19102, W17861, W19111);
not G20500 (W19103, W19562);
not G20501 (W19104, W19562);
nand G20502 (W19105, W19111, W19563);
not G20503 (W19106, W19108);
nand G20504 (W19107, W15842, W17197);
not G20505 (W19108, W19564);
nand G20506 (W19109, W18589, W19111);
not G20507 (W19110, W19112);
not G20508 (W19111, W18590);
not G20509 (W19112, W19565);
nor G20510 (W19113, W15842, W17861, W17197);
not G20511 (W19114, W19116);
nor G20512 (W19115, W15842, W19111);
not G20513 (W19116, W19566);
nor G20514 (W19117, W13464, W15763);
and G20515 (W19118, W11348, W11340);
nor G20516 (W19119, W19567, W19568, W19569);
nor G20517 (W19120, W19570, W19571, W19572);
nor G20518 (W19121, W19573, W19574, W19575);
and G20519 (W19122, W19576, W19577, W19578);
nor G20520 (W19123, W19579, W19580, W19581);
nor G20521 (W19124, W19582, W19583, W19584);
nor G20522 (W19125, W19585, W19586);
and G20523 (W19126, W19587, W19588, W19589);
and G20524 (W19127, W18597, I1561);
and G20525 (W19128, W19590, I1562);
and G20526 (W19129, W18597, W19591);
and G20527 (W19130, W19590, I1563);
and G20528 (W19131, W18597, I1564);
and G20529 (W19132, W19590, I1565);
nand G20530 (W19133, W19592, W19593);
or G20531 (W19134, W19594, W19595);
and G20532 (W19135, W19596, W19597);
and G20533 (W19136, W19598, W19599);
and G20534 (W19137, W19600, W19601);
and G20535 (W19138, W19602, I1566);
and G20536 (W19139, W19603, I1567);
and G20537 (W19140, W19604, W19605);
and G20538 (W19141, W19606, W19607);
and G20539 (W19142, W19590, I1568);
and G20540 (W19143, W18597, W19608);
nor G20541 (W19144, W19609, W19610);
nor G20542 (W19145, W19611, W19612, W19613);
nor G20543 (W19146, W19614, W19615, W19616);
and G20544 (W19147, W19617, W19618);
and G20545 (W19148, W19619, W17262);
and G20546 (W19149, W18597, W19620);
and G20547 (W19150, W19602, I1518);
and G20548 (W19151, W19603, I1569);
not G20549 (W19152, W19621);
not G20550 (W19153, W19622);
not G20551 (W19154, W19623);
not G20552 (W19155, W19624);
not G20553 (W19156, W19625);
not G20554 (W19157, W19626);
not G20555 (W19158, W5252);
not G20556 (W19159, W19627);
not G20557 (W19160, W19628);
not G20558 (W19161, W19629);
not G20559 (W19162, W19630);
not G20560 (W19163, W19631);
and G20561 (W19164, W18616, W19158, W18606);
and G20562 (W19165, W5252, W18621, W18610);
and G20563 (W19166, W19158, W18621, W18606);
not G20564 (W19167, W19632);
not G20565 (W19168, W19633);
not G20566 (W19169, W19634);
not G20567 (W19170, W4977);
not G20568 (W19171, W19635);
not G20569 (W19172, W19636);
not G20570 (W19173, W19637);
not G20571 (W19174, W19638);
not G20572 (W19175, W19639);
and G20573 (W19176, W18642, W19170, W18632);
and G20574 (W19177, W4977, W18647, W18636);
and G20575 (W19178, W19170, W18647, W18632);
not G20576 (W19179, W19640);
not G20577 (W19180, W19641);
not G20578 (W19181, W19642);
not G20579 (W19182, W4702);
not G20580 (W19183, W19643);
not G20581 (W19184, W19644);
not G20582 (W19185, W19645);
not G20583 (W19186, W19646);
not G20584 (W19187, W19647);
and G20585 (W19188, W18668, W19182, W18658);
and G20586 (W19189, W4702, W18673, W18662);
and G20587 (W19190, W19182, W18673, W18658);
not G20588 (W19191, W19648);
not G20589 (W19192, W19649);
not G20590 (W19193, W19650);
not G20591 (W19194, W4427);
not G20592 (W19195, W19651);
not G20593 (W19196, W19652);
not G20594 (W19197, W19653);
not G20595 (W19198, W19654);
not G20596 (W19199, W19655);
and G20597 (W19200, W18694, W19194, W18684);
and G20598 (W19201, W4427, W18699, W18688);
and G20599 (W19202, W19194, W18699, W18684);
nor G20600 (W19203, W19656, W19657, W19658);
not G20601 (W19204, W17327);
and G20602 (W19205, W19659, W17991, W17993);
and G20603 (W19206, W19660, W19661, W19662);
and G20604 (W19207, W15138, W8495);
and G20605 (W19208, W8544, W8492);
and G20606 (W19209, W13643, W8489);
and G20607 (W19210, W15138, W8486);
and G20608 (W19211, W8544, W8483);
and G20609 (W19212, W13643, W8480);
and G20610 (W19213, W15138, W8477);
and G20611 (W19214, W8544, W8474);
and G20612 (W19215, W13643, W8471);
and G20613 (W19216, W15138, W8540);
and G20614 (W19217, W8544, W8537);
and G20615 (W19218, W13643, W8534);
and G20616 (W19219, W15138, W8531);
and G20617 (W19220, W8544, W8528);
and G20618 (W19221, W13643, W8525);
and G20619 (W19222, W15138, W8522);
and G20620 (W19223, W8544, W8519);
and G20621 (W19224, W13643, W8516);
and G20622 (W19225, W13950, W9055);
and G20623 (W19226, W13951, W9052);
and G20624 (W19227, W9107, W9011);
and G20625 (W19228, W13950, W9061);
and G20626 (W19229, W13951, W9058);
and G20627 (W19230, W9107, W9015);
nor G20628 (W19231, W19663, W19664, W19665);
nor G20629 (W19232, W19666, W19667, W19668);
nor G20630 (W19233, W19669, W19670, W19671);
and G20631 (W19234, W13950, W9088);
and G20632 (W19235, W13951, W9082);
and G20633 (W19236, W9107, W9031);
and G20634 (W19237, W13950, W9100);
and G20635 (W19238, W13951, W9091);
and G20636 (W19239, W9107, W9039);
nor G20637 (W19240, W19672, W19673, W19674);
nor G20638 (W19241, W19675, W19676, W19677);
nor G20639 (W19242, W19678, W19679, W19680);
nor G20640 (W19243, W19681, W19682);
nor G20641 (W19244, W19683, W19684);
nor G20642 (W19245, W19685, W19686);
not G20643 (W19246, W19248);
and G20644 (W19247, W16647, W16676, W16705, W19687);
not G20645 (W19248, W19688);
nor G20646 (W19249, W19689, W19690, W19691);
nor G20647 (W19250, W19692, W19693);
and G20648 (W19251, W16672, W19694);
and G20649 (W19252, W16674, W19695);
and G20650 (W19253, W16682, W19696);
and G20651 (W19254, W16684, W19697);
and G20652 (W19255, W16688, W19698);
and G20653 (W19256, W16690, W19699);
and G20654 (W19257, W16638, W19700);
and G20655 (W19258, W16640, W19701);
and G20656 (W19259, W16645, W19702);
and G20657 (W19260, W16647, W19703);
nor G20658 (W19261, W19704, W19705);
not G20659 (W19262, W19264);
nand G20660 (W19263, W15195, W13982, W19706, W19707);
not G20661 (W19264, W19708);
and G20662 (W19265, W19707, W19709);
and G20663 (W19266, W19710, W19711);
and G20664 (W19267, W19712, W19713);
and G20665 (W19268, W19714, W19715);
not G20666 (W19269, W13983);
nand G20667 (W19270, W19716, W19717);
or G20668 (W19271, W19276, W19718);
or G20669 (W19272, W19273, W19719);
nand G20670 (W19273, W19720, W19721);
or G20671 (W19274, W19718, W19270);
or G20672 (W19275, W19276, W19719);
nand G20673 (W19276, W19722, W19723);
or G20674 (W19277, W19718, W19273);
or G20675 (W19278, W19719, W19270);
nand G20676 (W19279, W19724, W19725);
or G20677 (W19280, W19285, W19726);
or G20678 (W19281, W19282, W19727);
nand G20679 (W19282, W19728, W19729);
or G20680 (W19283, W19726, W19279);
or G20681 (W19284, W19285, W19727);
nand G20682 (W19285, W19730, W19731);
or G20683 (W19286, W19726, W19282);
or G20684 (W19287, W19727, W19279);
nor G20685 (W19288, W19732, W19733);
not G20686 (W19289, W19734);
or G20687 (W19290, W15274, W17422);
not G20688 (W19291, W4560);
not G20689 (W19292, W4560);
not G20690 (W19293, W4560);
nor G20691 (W19294, W19735, W19736, W19737);
not G20692 (W19295, W17473);
and G20693 (W19296, W19738, W18150, W18152);
and G20694 (W19297, W19739, W19740, W19741);
and G20695 (W19298, W15335, W9268);
and G20696 (W19299, W9317, W9265);
and G20697 (W19300, W13642, W9262);
and G20698 (W19301, W15335, W9259);
and G20699 (W19302, W9317, W9256);
and G20700 (W19303, W13642, W9253);
and G20701 (W19304, W15335, W9250);
and G20702 (W19305, W9317, W9247);
and G20703 (W19306, W13642, W9244);
and G20704 (W19307, W15335, W9313);
and G20705 (W19308, W9317, W9310);
and G20706 (W19309, W13642, W9307);
and G20707 (W19310, W15335, W9304);
and G20708 (W19311, W9317, W9301);
and G20709 (W19312, W13642, W9298);
and G20710 (W19313, W15335, W9295);
and G20711 (W19314, W9317, W9292);
and G20712 (W19315, W13642, W9289);
and G20713 (W19316, W14244, W9828);
and G20714 (W19317, W14245, W9825);
and G20715 (W19318, W9880, W9784);
and G20716 (W19319, W14244, W9834);
and G20717 (W19320, W14245, W9831);
and G20718 (W19321, W9880, W9788);
nor G20719 (W19322, W19742, W19743, W19744);
nor G20720 (W19323, W19745, W19746, W19747);
nor G20721 (W19324, W19748, W19749, W19750);
and G20722 (W19325, W14244, W9861);
and G20723 (W19326, W14245, W9855);
and G20724 (W19327, W9880, W9804);
and G20725 (W19328, W14244, W9873);
and G20726 (W19329, W14245, W9864);
and G20727 (W19330, W9880, W9812);
nor G20728 (W19331, W19751, W19752, W19753);
nor G20729 (W19332, W19754, W19755, W19756);
nor G20730 (W19333, W19757, W19758, W19759);
nor G20731 (W19334, W19760, W19761);
nor G20732 (W19335, W19762, W19763);
nor G20733 (W19336, W19764, W19765);
not G20734 (W19337, W19339);
and G20735 (W19338, W16802, W16831, W16860, W19766);
not G20736 (W19339, W19767);
nor G20737 (W19340, W19768, W19769, W19770);
nor G20738 (W19341, W19771, W19772);
and G20739 (W19342, W16827, W19773);
and G20740 (W19343, W16829, W19774);
and G20741 (W19344, W16837, W19775);
and G20742 (W19345, W16839, W19776);
and G20743 (W19346, W16843, W19777);
and G20744 (W19347, W16845, W19778);
and G20745 (W19348, W16793, W19779);
and G20746 (W19349, W16795, W19780);
and G20747 (W19350, W16800, W19781);
and G20748 (W19351, W16802, W19782);
nor G20749 (W19352, W19783, W19784);
not G20750 (W19353, W19355);
nand G20751 (W19354, W15389, W14276, W19785, W19786);
not G20752 (W19355, W19787);
and G20753 (W19356, W19786, W19788);
and G20754 (W19357, W19789, W19790);
and G20755 (W19358, W19791, W19792);
and G20756 (W19359, W19793, W19794);
not G20757 (W19360, W14277);
nand G20758 (W19361, W19795, W19796);
or G20759 (W19362, W19367, W19797);
or G20760 (W19363, W19364, W19798);
nand G20761 (W19364, W19799, W19800);
or G20762 (W19365, W19797, W19361);
or G20763 (W19366, W19367, W19798);
nand G20764 (W19367, W19801, W19802);
or G20765 (W19368, W19797, W19364);
or G20766 (W19369, W19798, W19361);
nand G20767 (W19370, W19803, W19804);
or G20768 (W19371, W19376, W19805);
or G20769 (W19372, W19373, W19806);
nand G20770 (W19373, W19807, W19808);
or G20771 (W19374, W19805, W19370);
or G20772 (W19375, W19376, W19806);
nand G20773 (W19376, W19809, W19810);
or G20774 (W19377, W19805, W19373);
or G20775 (W19378, W19806, W19370);
nor G20776 (W19379, W19811, W19812);
not G20777 (W19380, W19813);
or G20778 (W19381, W15467, W17568);
not G20779 (W19382, W4835);
not G20780 (W19383, W4835);
not G20781 (W19384, W4835);
nor G20782 (W19385, W19814, W19815, W19816);
not G20783 (W19386, W17619);
and G20784 (W19387, W19817, W18309, W18311);
and G20785 (W19388, W19818, W19819, W19820);
and G20786 (W19389, W15528, W10041);
and G20787 (W19390, W10090, W10038);
and G20788 (W19391, W13641, W10035);
and G20789 (W19392, W15528, W10032);
and G20790 (W19393, W10090, W10029);
and G20791 (W19394, W13641, W10026);
and G20792 (W19395, W15528, W10023);
and G20793 (W19396, W10090, W10020);
and G20794 (W19397, W13641, W10017);
and G20795 (W19398, W15528, W10086);
and G20796 (W19399, W10090, W10083);
and G20797 (W19400, W13641, W10080);
and G20798 (W19401, W15528, W10077);
and G20799 (W19402, W10090, W10074);
and G20800 (W19403, W13641, W10071);
and G20801 (W19404, W15528, W10068);
and G20802 (W19405, W10090, W10065);
and G20803 (W19406, W13641, W10062);
and G20804 (W19407, W14537, W10598);
and G20805 (W19408, W14538, W10595);
and G20806 (W19409, W10653, W10553);
and G20807 (W19410, W14537, W10604);
and G20808 (W19411, W14538, W10601);
and G20809 (W19412, W10653, W10557);
nor G20810 (W19413, W19821, W19822, W19823);
nor G20811 (W19414, W19824, W19825, W19826);
nor G20812 (W19415, W19827, W19828, W19829);
and G20813 (W19416, W14537, W10631);
and G20814 (W19417, W14538, W10625);
and G20815 (W19418, W10653, W10573);
and G20816 (W19419, W14537, W10643);
and G20817 (W19420, W14538, W10634);
and G20818 (W19421, W10653, W10581);
nor G20819 (W19422, W19830, W19831, W19832);
nor G20820 (W19423, W19833, W19834, W19835);
nor G20821 (W19424, W19836, W19837, W19838);
nor G20822 (W19425, W19839, W19840);
nor G20823 (W19426, W19841, W19842);
nor G20824 (W19427, W19843, W19844);
not G20825 (W19428, W19430);
and G20826 (W19429, W16957, W16986, W17015, W19845);
not G20827 (W19430, W19846);
nor G20828 (W19431, W19847, W19848, W19849);
nor G20829 (W19432, W19850, W19851);
and G20830 (W19433, W16982, W19852);
and G20831 (W19434, W16984, W19853);
and G20832 (W19435, W16992, W19854);
and G20833 (W19436, W16994, W19855);
and G20834 (W19437, W16998, W19856);
and G20835 (W19438, W17000, W19857);
and G20836 (W19439, W16948, W19858);
and G20837 (W19440, W16950, W19859);
and G20838 (W19441, W16955, W19860);
and G20839 (W19442, W16957, W19861);
nor G20840 (W19443, W19862, W19863);
not G20841 (W19444, W19446);
nand G20842 (W19445, W15582, W14569, W19864, W19865);
not G20843 (W19446, W19866);
and G20844 (W19447, W19865, W19867);
and G20845 (W19448, W19868, W19869);
and G20846 (W19449, W19870, W19871);
and G20847 (W19450, W19872, W19873);
not G20848 (W19451, W14570);
nand G20849 (W19452, W19874, W19875);
or G20850 (W19453, W19458, W19876);
or G20851 (W19454, W19455, W19877);
nand G20852 (W19455, W19878, W19879);
or G20853 (W19456, W19876, W19452);
or G20854 (W19457, W19458, W19877);
nand G20855 (W19458, W19880, W19881);
or G20856 (W19459, W19876, W19455);
or G20857 (W19460, W19877, W19452);
nand G20858 (W19461, W19882, W19883);
or G20859 (W19462, W19467, W19884);
or G20860 (W19463, W19464, W19885);
nand G20861 (W19464, W19886, W19887);
or G20862 (W19465, W19884, W19461);
or G20863 (W19466, W19467, W19885);
nand G20864 (W19467, W19888, W19889);
or G20865 (W19468, W19884, W19464);
or G20866 (W19469, W19885, W19461);
nor G20867 (W19470, W19890, W19891);
not G20868 (W19471, W19892);
or G20869 (W19472, W15660, W17714);
not G20870 (W19473, W5110);
not G20871 (W19474, W5110);
not G20872 (W19475, W5110);
nor G20873 (W19476, W19893, W19894, W19895);
not G20874 (W19477, W17766);
and G20875 (W19478, W19896, W18469, W18471);
and G20876 (W19479, W19897, W19898, W19899);
and G20877 (W19480, W15721, W10814);
and G20878 (W19481, W10863, W10811);
and G20879 (W19482, W13640, W10808);
and G20880 (W19483, W15721, W10805);
and G20881 (W19484, W10863, W10802);
and G20882 (W19485, W13640, W10799);
and G20883 (W19486, W15721, W10796);
and G20884 (W19487, W10863, W10793);
and G20885 (W19488, W13640, W10790);
and G20886 (W19489, W15721, W10859);
and G20887 (W19490, W10863, W10856);
and G20888 (W19491, W13640, W10853);
and G20889 (W19492, W15721, W10850);
and G20890 (W19493, W10863, W10847);
and G20891 (W19494, W13640, W10844);
and G20892 (W19495, W15721, W10841);
and G20893 (W19496, W10863, W10838);
and G20894 (W19497, W13640, W10835);
and G20895 (W19498, W14808, W11368);
and G20896 (W19499, W14809, W11365);
and G20897 (W19500, W11426, W11422);
and G20898 (W19501, W14808, W11374);
and G20899 (W19502, W14809, W11371);
and G20900 (W19503, W11426, W11326);
nor G20901 (W19504, W19900, W19901, W19902);
nor G20902 (W19505, W19903, W19904, W19905);
nor G20903 (W19506, W19906, W19907, W19908);
and G20904 (W19507, W14808, W11401);
and G20905 (W19508, W14809, W11395);
and G20906 (W19509, W11426, W11342);
and G20907 (W19510, W14808, W11413);
and G20908 (W19511, W14809, W11404);
and G20909 (W19512, W11426, W11350);
nor G20910 (W19513, W19909, W19910, W19911);
nor G20911 (W19514, W19912, W19913, W19914);
nor G20912 (W19515, W19915, W19916, W19917);
nor G20913 (W19516, W19918, W19919);
nor G20914 (W19517, W19920, W19921);
nor G20915 (W19518, W19922, W19923);
not G20916 (W19519, W19521);
and G20917 (W19520, W17112, W17141, W17170, W19924);
not G20918 (W19521, W19925);
nor G20919 (W19522, W19926, W19927, W19928);
nor G20920 (W19523, W19929, W19930);
and G20921 (W19524, W17137, W19931);
and G20922 (W19525, W17139, W19932);
and G20923 (W19526, W17147, W19933);
and G20924 (W19527, W17149, W19934);
and G20925 (W19528, W17153, W19935);
and G20926 (W19529, W17155, W19936);
and G20927 (W19530, W17103, W19937);
and G20928 (W19531, W17105, W19938);
and G20929 (W19532, W17110, W19939);
and G20930 (W19533, W17112, W19940);
nor G20931 (W19534, W19941, W19942);
not G20932 (W19535, W19537);
nand G20933 (W19536, W15764, W14840, W19943, W19944);
not G20934 (W19537, W19945);
and G20935 (W19538, W19944, W19946);
and G20936 (W19539, W19947, W19948);
and G20937 (W19540, W19949, W19950);
and G20938 (W19541, W19951, W19952);
not G20939 (W19542, W14841);
nand G20940 (W19543, W19953, W19954);
or G20941 (W19544, W19549, W19955);
or G20942 (W19545, W19546, W19956);
nand G20943 (W19546, W19957, W19958);
or G20944 (W19547, W19955, W19543);
or G20945 (W19548, W19549, W19956);
nand G20946 (W19549, W19959, W19960);
or G20947 (W19550, W19955, W19546);
or G20948 (W19551, W19956, W19543);
nand G20949 (W19552, W19961, W19962);
or G20950 (W19553, W19558, W19963);
or G20951 (W19554, W19555, W19964);
nand G20952 (W19555, W19965, W19966);
or G20953 (W19556, W19963, W19552);
or G20954 (W19557, W19558, W19964);
nand G20955 (W19558, W19967, W19968);
or G20956 (W19559, W19963, W19555);
or G20957 (W19560, W19964, W19552);
nor G20958 (W19561, W19969, W19970);
not G20959 (W19562, W19971);
or G20960 (W19563, W15842, W17861);
not G20961 (W19564, W5385);
not G20962 (W19565, W5385);
not G20963 (W19566, W5385);
and G20964 (W19567, W19596, W19972);
and G20965 (W19568, W19598, W19973);
and G20966 (W19569, W19600, W19974);
and G20967 (W19570, W19602, I1393);
and G20968 (W19571, W19603, I1570);
and G20969 (W19572, W19604, W19975);
and G20970 (W19573, W19606, W19976);
and G20971 (W19574, W19590, I1571);
and G20972 (W19575, W18597, I1572);
nor G20973 (W19576, W19977, W19978);
nor G20974 (W19577, W19979, W19980, W19981);
nor G20975 (W19578, W19982, W19983, W19984);
and G20976 (W19579, W19598, I1221);
and G20977 (W19580, W19600, I1018);
and G20978 (W19581, W19985, I1019);
and G20979 (W19582, W19602, I1573);
and G20980 (W19583, W19604, I1219);
and G20981 (W19584, W19596, I1220);
and G20982 (W19585, W19590, I1574);
and G20983 (W19586, W18597, I1575);
nand G20984 (W19587, I618, W19986);
nor G20985 (W19588, W19987, W19988, W19989);
nor G20986 (W19589, W19990, W19991, W19992);
not G20987 (W19590, W19993);
not G20988 (W19591, I1576);
nor G20989 (W19592, W19994, W19995, W19996, W19997);
not G20990 (W19593, W19998);
not G20991 (W19594, W19999);
not G20992 (W19595, W20000);
not G20993 (W19596, W20001);
not G20994 (W19597, W10956);
not G20995 (W19598, W20002);
not G20996 (W19599, W10959);
not G20997 (W19600, W20003);
not G20998 (W19601, W10179);
not G20999 (W19602, W20004);
not G21000 (W19603, W20005);
not G21001 (W19604, W20006);
not G21002 (W19605, W10952);
not G21003 (W19606, W20007);
not G21004 (W19607, W20008);
not G21005 (W19608, I1577);
and G21006 (W19609, W20009, W20010);
and G21007 (W19610, W19986, W20011);
and G21008 (W19611, W20012, W20013);
and G21009 (W19612, W20014, W20015);
and G21010 (W19613, W20016, W20017);
and G21011 (W19614, W19985, W20018);
and G21012 (W19615, W20019, W20020);
and G21013 (W19616, W20021, W20022);
not G21014 (W19617, W20023);
not G21015 (W19618, W20024);
not G21016 (W19619, W20025);
not G21017 (W19620, I1578);
nand G21018 (W19621, W20026, W19593);
nand G21019 (W19622, W20027, W19593);
not G21020 (W19623, W19606);
nor G21021 (W19624, W20028, W20029, W20030);
not G21022 (W19625, W19630);
not G21023 (W19626, W19629);
not G21024 (W19627, W19624);
not G21025 (W19628, W19631);
nor G21026 (W19629, W20031, W20032, W20033);
nor G21027 (W19630, W20034, W20035, W20036);
nor G21028 (W19631, W20037, W20038, W20039);
nor G21029 (W19632, W20040, W20041, W20042);
not G21030 (W19633, W19638);
not G21031 (W19634, W19637);
not G21032 (W19635, W19632);
not G21033 (W19636, W19639);
nor G21034 (W19637, W20043, W20044, W20045);
nor G21035 (W19638, W20046, W20047, W20048);
nor G21036 (W19639, W20049, W20050, W20051);
nor G21037 (W19640, W20052, W20053, W20054);
not G21038 (W19641, W19646);
not G21039 (W19642, W19645);
not G21040 (W19643, W19640);
not G21041 (W19644, W19647);
nor G21042 (W19645, W20055, W20056, W20057);
nor G21043 (W19646, W20058, W20059, W20060);
nor G21044 (W19647, W20061, W20062, W20063);
nor G21045 (W19648, W20064, W20065, W20066);
not G21046 (W19649, W19654);
not G21047 (W19650, W19653);
not G21048 (W19651, W19648);
not G21049 (W19652, W19655);
nor G21050 (W19653, W20067, W20068, W20069);
nor G21051 (W19654, W20070, W20071, W20072);
nor G21052 (W19655, W20073, W20074, W20075);
and G21053 (W19656, W15138, W8420);
and G21054 (W19657, W8544, W8417);
and G21055 (W19658, W13643, W8414);
not G21056 (W19659, W17989);
not G21057 (W19660, W17981);
not G21058 (W19661, W17983);
not G21059 (W19662, W17985);
and G21060 (W19663, W13950, W9094);
and G21061 (W19664, W13951, W9085);
and G21062 (W19665, W9107, W9035);
and G21063 (W19666, W13950, W9103);
and G21064 (W19667, W13951, W9097);
and G21065 (W19668, W9107, W9043);
and G21066 (W19669, W13950, W9049);
and G21067 (W19670, W13951, W9046);
and G21068 (W19671, W9107, W9007);
and G21069 (W19672, W13950, W9067);
and G21070 (W19673, W13951, W9064);
and G21071 (W19674, W9107, W9019);
and G21072 (W19675, W13950, W9073);
and G21073 (W19676, W13951, W9070);
and G21074 (W19677, W9107, W9023);
and G21075 (W19678, W13950, W9079);
and G21076 (W19679, W13951, W9076);
and G21077 (W19680, W9107, W9027);
and G21078 (W19681, W16666, W20076);
and G21079 (W19682, W16664, W20077);
and G21080 (W19683, W16652, W20078);
and G21081 (W19684, W16654, W20079);
and G21082 (W19685, W16660, W20080);
and G21083 (W19686, W16658, W20081);
and G21084 (W19687, W16654, W16684, W16658);
not G21085 (W19688, W17356);
and G21086 (W19689, W12210, W8886);
and G21087 (W19690, W12211, W8883);
and G21088 (W19691, W12212, W8880);
and G21089 (W19692, W16670, W20082);
and G21090 (W19693, W16668, W20083);
not G21091 (W19694, W19695);
not G21092 (W19695, W20084);
not G21093 (W19696, W19697);
not G21094 (W19697, W20085);
not G21095 (W19698, W19699);
not G21096 (W19699, W20086);
not G21097 (W19700, W19701);
not G21098 (W19701, W20087);
not G21099 (W19702, W19703);
not G21100 (W19703, W20088);
and G21101 (W19704, W20089, W20090);
and G21102 (W19705, W20091, W20092);
not G21103 (W19706, W18765);
not G21104 (W19707, W18766);
not G21105 (W19708, W13983);
not G21106 (W19709, W19711);
nor G21107 (W19710, W18766, W20093);
not G21108 (W19711, W20094);
nor G21109 (W19712, W17422, W20095);
not G21110 (W19713, W19715);
nor G21111 (W19714, W18765, W20091, W20096);
not G21112 (W19715, W20097);
nand G21113 (W19716, W16672, W20098);
nand G21114 (W19717, W9033, W20098);
nand G21115 (W19718, W20099, W20100);
nand G21116 (W19719, W20101, W20102);
nand G21117 (W19720, W16690, W20103);
nand G21118 (W19721, W9013, W20103);
nand G21119 (W19722, W16647, W20104);
nand G21120 (W19723, W9029, W20104);
nand G21121 (W19724, W16654, W20105);
nand G21122 (W19725, W9041, W20105);
nand G21123 (W19726, W20106, W20107);
nand G21124 (W19727, W20108, W20109);
nand G21125 (W19728, W16664, W20110);
nand G21126 (W19729, W9017, W20110);
nand G21127 (W19730, W16676, W20111);
nand G21128 (W19731, W9037, W20111);
or G21129 (W19732, W19718, W19276, W20112);
or G21130 (W19733, W19726, W19285, W20113);
not G21131 (W19734, W4560);
and G21132 (W19735, W15335, W9193);
and G21133 (W19736, W9317, W9190);
and G21134 (W19737, W13642, W9187);
not G21135 (W19738, W18148);
not G21136 (W19739, W18140);
not G21137 (W19740, W18142);
not G21138 (W19741, W18144);
and G21139 (W19742, W14244, W9867);
and G21140 (W19743, W14245, W9858);
and G21141 (W19744, W9880, W9808);
and G21142 (W19745, W14244, W9876);
and G21143 (W19746, W14245, W9870);
and G21144 (W19747, W9880, W9816);
and G21145 (W19748, W14244, W9822);
and G21146 (W19749, W14245, W9819);
and G21147 (W19750, W9880, W9780);
and G21148 (W19751, W14244, W9840);
and G21149 (W19752, W14245, W9837);
and G21150 (W19753, W9880, W9792);
and G21151 (W19754, W14244, W9846);
and G21152 (W19755, W14245, W9843);
and G21153 (W19756, W9880, W9796);
and G21154 (W19757, W14244, W9852);
and G21155 (W19758, W14245, W9849);
and G21156 (W19759, W9880, W9800);
and G21157 (W19760, W16821, W20114);
and G21158 (W19761, W16819, W20115);
and G21159 (W19762, W16807, W20116);
and G21160 (W19763, W16809, W20117);
and G21161 (W19764, W16815, W20118);
and G21162 (W19765, W16813, W20119);
and G21163 (W19766, W16809, W16839, W16813);
not G21164 (W19767, W17502);
and G21165 (W19768, W12616, W9659);
and G21166 (W19769, W12617, W9656);
and G21167 (W19770, W12618, W9653);
and G21168 (W19771, W16825, W20120);
and G21169 (W19772, W16823, W20121);
not G21170 (W19773, W19774);
not G21171 (W19774, W20122);
not G21172 (W19775, W19776);
not G21173 (W19776, W20123);
not G21174 (W19777, W19778);
not G21175 (W19778, W20124);
not G21176 (W19779, W19780);
not G21177 (W19780, W20125);
not G21178 (W19781, W19782);
not G21179 (W19782, W20126);
and G21180 (W19783, W20127, W20128);
and G21181 (W19784, W20129, W20130);
not G21182 (W19785, W18867);
not G21183 (W19786, W18868);
not G21184 (W19787, W14277);
not G21185 (W19788, W19790);
nor G21186 (W19789, W18868, W20131);
not G21187 (W19790, W20132);
nor G21188 (W19791, W17568, W20133);
not G21189 (W19792, W19794);
nor G21190 (W19793, W18867, W20129, W20134);
not G21191 (W19794, W20135);
nand G21192 (W19795, W16827, W20136);
nand G21193 (W19796, W9806, W20136);
nand G21194 (W19797, W20137, W20138);
nand G21195 (W19798, W20139, W20140);
nand G21196 (W19799, W16845, W20141);
nand G21197 (W19800, W9786, W20141);
nand G21198 (W19801, W16802, W20142);
nand G21199 (W19802, W9802, W20142);
nand G21200 (W19803, W16809, W20143);
nand G21201 (W19804, W9814, W20143);
nand G21202 (W19805, W20144, W20145);
nand G21203 (W19806, W20146, W20147);
nand G21204 (W19807, W16819, W20148);
nand G21205 (W19808, W9790, W20148);
nand G21206 (W19809, W16831, W20149);
nand G21207 (W19810, W9810, W20149);
or G21208 (W19811, W19797, W19367, W20150);
or G21209 (W19812, W19805, W19376, W20151);
not G21210 (W19813, W4835);
and G21211 (W19814, W15528, W9966);
and G21212 (W19815, W10090, W9963);
and G21213 (W19816, W13641, W9960);
not G21214 (W19817, W18307);
not G21215 (W19818, W18299);
not G21216 (W19819, W18301);
not G21217 (W19820, W18303);
and G21218 (W19821, W14537, W10637);
and G21219 (W19822, W14538, W10628);
and G21220 (W19823, W10653, W10577);
and G21221 (W19824, W14537, W10646);
and G21222 (W19825, W14538, W10640);
and G21223 (W19826, W10653, W10585);
and G21224 (W19827, W14537, W10592);
and G21225 (W19828, W14538, W10589);
and G21226 (W19829, W10653, W10649);
and G21227 (W19830, W14537, W10610);
and G21228 (W19831, W14538, W10607);
and G21229 (W19832, W10653, W10561);
and G21230 (W19833, W14537, W10616);
and G21231 (W19834, W14538, W10613);
and G21232 (W19835, W10653, W10565);
and G21233 (W19836, W14537, W10622);
and G21234 (W19837, W14538, W10619);
and G21235 (W19838, W10653, W10569);
and G21236 (W19839, W16976, W20152);
and G21237 (W19840, W16974, W20153);
and G21238 (W19841, W16962, W20154);
and G21239 (W19842, W16964, W20155);
and G21240 (W19843, W16970, W20156);
and G21241 (W19844, W16968, W20157);
and G21242 (W19845, W16964, W16994, W16968);
not G21243 (W19846, W17648);
and G21244 (W19847, W13022, W10432);
and G21245 (W19848, W13023, W10429);
and G21246 (W19849, W13024, W10426);
and G21247 (W19850, W16980, W20158);
and G21248 (W19851, W16978, W20159);
not G21249 (W19852, W19853);
not G21250 (W19853, W20160);
not G21251 (W19854, W19855);
not G21252 (W19855, W20161);
not G21253 (W19856, W19857);
not G21254 (W19857, W20162);
not G21255 (W19858, W19859);
not G21256 (W19859, W20163);
not G21257 (W19860, W19861);
not G21258 (W19861, W20164);
and G21259 (W19862, W20165, W20166);
and G21260 (W19863, W20167, W20168);
not G21261 (W19864, W18969);
not G21262 (W19865, W18970);
not G21263 (W19866, W14570);
not G21264 (W19867, W19869);
nor G21265 (W19868, W18970, W20169);
not G21266 (W19869, W20170);
nor G21267 (W19870, W17714, W20171);
not G21268 (W19871, W19873);
nor G21269 (W19872, W18969, W20167, W20172);
not G21270 (W19873, W20173);
nand G21271 (W19874, W16982, W20174);
nand G21272 (W19875, W10575, W20174);
nand G21273 (W19876, W20175, W20176);
nand G21274 (W19877, W20177, W20178);
nand G21275 (W19878, W17000, W20179);
nand G21276 (W19879, W10555, W20179);
nand G21277 (W19880, W16957, W20180);
nand G21278 (W19881, W10571, W20180);
nand G21279 (W19882, W16964, W20181);
nand G21280 (W19883, W10583, W20181);
nand G21281 (W19884, W20182, W20183);
nand G21282 (W19885, W20184, W20185);
nand G21283 (W19886, W16974, W20186);
nand G21284 (W19887, W10559, W20186);
nand G21285 (W19888, W16986, W20187);
nand G21286 (W19889, W10579, W20187);
or G21287 (W19890, W19876, W19458, W20188);
or G21288 (W19891, W19884, W19467, W20189);
not G21289 (W19892, W5110);
and G21290 (W19893, W15721, W10739);
and G21291 (W19894, W10863, W10736);
and G21292 (W19895, W13640, W10733);
not G21293 (W19896, W18467);
not G21294 (W19897, W18459);
not G21295 (W19898, W18461);
not G21296 (W19899, W18463);
and G21297 (W19900, W14808, W11407);
and G21298 (W19901, W14809, W11398);
and G21299 (W19902, W11426, W11346);
and G21300 (W19903, W14808, W11416);
and G21301 (W19904, W14809, W11410);
and G21302 (W19905, W11426, W11354);
and G21303 (W19906, W14808, W11361);
and G21304 (W19907, W14809, W11358);
and G21305 (W19908, W11426, W11419);
and G21306 (W19909, W14808, W11380);
and G21307 (W19910, W14809, W11377);
and G21308 (W19911, W11426, W11330);
and G21309 (W19912, W14808, W11386);
and G21310 (W19913, W14809, W11383);
and G21311 (W19914, W11426, W11334);
and G21312 (W19915, W14808, W11392);
and G21313 (W19916, W14809, W11389);
and G21314 (W19917, W11426, W11338);
and G21315 (W19918, W17131, W20190);
and G21316 (W19919, W17129, W20191);
and G21317 (W19920, W17117, W20192);
and G21318 (W19921, W17119, W20193);
and G21319 (W19922, W17125, W20194);
and G21320 (W19923, W17123, W20195);
and G21321 (W19924, W17119, W17149, W17123);
not G21322 (W19925, W17795);
and G21323 (W19926, W13417, W11205);
and G21324 (W19927, W13418, W11202);
and G21325 (W19928, W13419, W11199);
and G21326 (W19929, W17135, W20196);
and G21327 (W19930, W17133, W20197);
not G21328 (W19931, W19932);
not G21329 (W19932, W20198);
not G21330 (W19933, W19934);
not G21331 (W19934, W20199);
not G21332 (W19935, W19936);
not G21333 (W19936, W20200);
not G21334 (W19937, W19938);
not G21335 (W19938, W20201);
not G21336 (W19939, W19940);
not G21337 (W19940, W20202);
and G21338 (W19941, W20203, W20204);
and G21339 (W19942, W20205, W20206);
not G21340 (W19943, W19071);
not G21341 (W19944, W19072);
not G21342 (W19945, W14841);
not G21343 (W19946, W19948);
nor G21344 (W19947, W19072, W20207);
not G21345 (W19948, W20208);
nor G21346 (W19949, W17861, W20209);
not G21347 (W19950, W19952);
nor G21348 (W19951, W19071, W20205, W20210);
not G21349 (W19952, W20211);
nand G21350 (W19953, W17137, W20212);
nand G21351 (W19954, W11344, W20212);
nand G21352 (W19955, W20213, W20214);
nand G21353 (W19956, W20215, W20216);
nand G21354 (W19957, W17155, W20217);
nand G21355 (W19958, W11324, W20217);
nand G21356 (W19959, W17112, W20218);
nand G21357 (W19960, W11340, W20218);
nand G21358 (W19961, W17119, W20219);
nand G21359 (W19962, W11352, W20219);
nand G21360 (W19963, W20220, W20221);
nand G21361 (W19964, W20222, W20223);
nand G21362 (W19965, W17129, W20224);
nand G21363 (W19966, W11328, W20224);
nand G21364 (W19967, W17141, W20225);
nand G21365 (W19968, W11348, W20225);
or G21366 (W19969, W19955, W19549, W20226);
or G21367 (W19970, W19963, W19558, W20227);
not G21368 (W19971, W5385);
not G21369 (W19972, W10932);
not G21370 (W19973, W10935);
not G21371 (W19974, W10155);
not G21372 (W19975, W10928);
not G21373 (W19976, W20228);
and G21374 (W19977, W20009, W20229);
and G21375 (W19978, W19986, W20230);
and G21376 (W19979, W20012, W20231);
and G21377 (W19980, W20014, W20232);
and G21378 (W19981, W20016, W20233);
and G21379 (W19982, W19985, W20234);
and G21380 (W19983, W20019, W20235);
and G21381 (W19984, W20021, W20236);
not G21382 (W19985, W20237);
not G21383 (W19986, W20238);
and G21384 (W19987, W20014, I819);
and G21385 (W19988, W20016, I616);
and G21386 (W19989, W20009, I617);
and G21387 (W19990, W20019, I1020);
and G21388 (W19991, W20021, I817);
and G21389 (W19992, W20012, I818);
nand G21390 (W19993, W20239, W19593);
not G21391 (W19994, W20240);
not G21392 (W19995, I1579);
not G21393 (W19996, W20241);
not G21394 (W19997, I1580);
nand G21395 (W19998, W20242, W20243, W20244, W20245);
not G21396 (W19999, W20246);
not G21397 (W20000, W20247);
nand G21398 (W20001, W20248, W20249);
nand G21399 (W20002, W20250, W20249);
nand G21400 (W20003, W20251, W20249);
nand G21401 (W20004, W20252, W19593);
nand G21402 (W20005, W20253, W19593);
nand G21403 (W20006, W20254, W20249);
nand G21404 (W20007, W20254, W19593);
not G21405 (W20008, W20255);
not G21406 (W20009, W20256);
not G21407 (W20010, W8637);
not G21408 (W20011, W8640);
not G21409 (W20012, W20257);
not G21410 (W20013, W9410);
not G21411 (W20014, W20258);
not G21412 (W20015, W9413);
not G21413 (W20016, W20259);
not G21414 (W20017, W8633);
not G21415 (W20018, W10183);
not G21416 (W20019, W20260);
not G21417 (W20020, W10186);
not G21418 (W20021, W20261);
not G21419 (W20022, W9406);
nand G21420 (W20023, W20252, W20249);
not G21421 (W20024, W20262);
nand G21422 (W20025, W20263, W20249);
nor G21423 (W20026, W19994, W20264, W19996, W19997);
nor G21424 (W20027, W20265, W20264, W19996, W19997);
and G21425 (W20028, I170, I1581);
and G21426 (W20029, I169, I1582);
and G21427 (W20030, I1583, I1584);
and G21428 (W20031, I170, I1585);
and G21429 (W20032, I169, I1586);
and G21430 (W20033, I1583, I1587);
and G21431 (W20034, I170, I1588);
and G21432 (W20035, I169, I1589);
and G21433 (W20036, I1583, I1590);
and G21434 (W20037, I170, I1591);
and G21435 (W20038, I169, I1592);
and G21436 (W20039, I1583, I1593);
and G21437 (W20040, I121, I1594);
and G21438 (W20041, I120, I1595);
and G21439 (W20042, I1596, I1597);
and G21440 (W20043, I121, I1598);
and G21441 (W20044, I120, I1599);
and G21442 (W20045, I1596, I1600);
and G21443 (W20046, I121, I1601);
and G21444 (W20047, I120, I1602);
and G21445 (W20048, I1596, I1603);
and G21446 (W20049, I121, I1604);
and G21447 (W20050, I120, I1605);
and G21448 (W20051, I1596, I1606);
and G21449 (W20052, I72, I1607);
and G21450 (W20053, I71, I1608);
and G21451 (W20054, I1609, I1610);
and G21452 (W20055, I72, I1611);
and G21453 (W20056, I71, I1612);
and G21454 (W20057, I1609, I1613);
and G21455 (W20058, I72, I1614);
and G21456 (W20059, I71, I1615);
and G21457 (W20060, I1609, I1616);
and G21458 (W20061, I72, I1617);
and G21459 (W20062, I71, I1618);
and G21460 (W20063, I1609, I1619);
and G21461 (W20064, I23, I1620);
and G21462 (W20065, I22, I1621);
and G21463 (W20066, I1622, I1623);
and G21464 (W20067, I23, I1624);
and G21465 (W20068, I22, I1625);
and G21466 (W20069, I1622, I1626);
and G21467 (W20070, I23, I1627);
and G21468 (W20071, I22, I1628);
and G21469 (W20072, I1622, I1629);
and G21470 (W20073, I23, I1630);
and G21471 (W20074, I22, I1631);
and G21472 (W20075, I1622, I1632);
not G21473 (W20076, W20077);
not G21474 (W20077, W20266);
not G21475 (W20078, W20079);
not G21476 (W20079, W20267);
not G21477 (W20080, W20081);
not G21478 (W20081, W20268);
not G21479 (W20082, W20083);
not G21480 (W20083, W20269);
not G21481 (W20084, W17356);
not G21482 (W20085, W17356);
not G21483 (W20086, W17356);
not G21484 (W20087, W17356);
not G21485 (W20088, W17356);
nand G21486 (W20089, W19706, W19707, W16702);
not G21487 (W20090, W20092);
or G21488 (W20091, W20270, W17422);
not G21489 (W20092, W20271);
and G21490 (W20093, W19706, W17390);
not G21491 (W20094, W13982);
and G21492 (W20095, W12099, W18757);
and G21493 (W20096, W17390, W15243, W18757);
not G21494 (W20097, W13982);
nand G21495 (W20098, W16672, W9033);
nand G21496 (W20099, W16640, W20272);
nand G21497 (W20100, W9021, W20272);
nand G21498 (W20101, W16684, W20273);
nand G21499 (W20102, W9005, W20273);
nand G21500 (W20103, W16690, W9013);
nand G21501 (W20104, W16647, W9029);
nand G21502 (W20105, W16654, W9041);
nand G21503 (W20106, W16668, W20274);
nand G21504 (W20107, W9025, W20274);
nand G21505 (W20108, W16658, W20275);
nand G21506 (W20109, W9009, W20275);
nand G21507 (W20110, W16664, W9017);
nand G21508 (W20111, W16676, W9037);
or G21509 (W20112, W19270, W19719, W19273);
or G21510 (W20113, W19279, W19727, W19282);
not G21511 (W20114, W20115);
not G21512 (W20115, W20276);
not G21513 (W20116, W20117);
not G21514 (W20117, W20277);
not G21515 (W20118, W20119);
not G21516 (W20119, W20278);
not G21517 (W20120, W20121);
not G21518 (W20121, W20279);
not G21519 (W20122, W17502);
not G21520 (W20123, W17502);
not G21521 (W20124, W17502);
not G21522 (W20125, W17502);
not G21523 (W20126, W17502);
nand G21524 (W20127, W19785, W19786, W16857);
not G21525 (W20128, W20130);
or G21526 (W20129, W20280, W17568);
not G21527 (W20130, W20281);
and G21528 (W20131, W19785, W17536);
not G21529 (W20132, W14276);
and G21530 (W20133, W12505, W18859);
and G21531 (W20134, W17536, W15437, W18859);
not G21532 (W20135, W14276);
nand G21533 (W20136, W16827, W9806);
nand G21534 (W20137, W16795, W20282);
nand G21535 (W20138, W9794, W20282);
nand G21536 (W20139, W16839, W20283);
nand G21537 (W20140, W9778, W20283);
nand G21538 (W20141, W16845, W9786);
nand G21539 (W20142, W16802, W9802);
nand G21540 (W20143, W16809, W9814);
nand G21541 (W20144, W16823, W20284);
nand G21542 (W20145, W9798, W20284);
nand G21543 (W20146, W16813, W20285);
nand G21544 (W20147, W9782, W20285);
nand G21545 (W20148, W16819, W9790);
nand G21546 (W20149, W16831, W9810);
or G21547 (W20150, W19361, W19798, W19364);
or G21548 (W20151, W19370, W19806, W19373);
not G21549 (W20152, W20153);
not G21550 (W20153, W20286);
not G21551 (W20154, W20155);
not G21552 (W20155, W20287);
not G21553 (W20156, W20157);
not G21554 (W20157, W20288);
not G21555 (W20158, W20159);
not G21556 (W20159, W20289);
not G21557 (W20160, W17648);
not G21558 (W20161, W17648);
not G21559 (W20162, W17648);
not G21560 (W20163, W17648);
not G21561 (W20164, W17648);
nand G21562 (W20165, W19864, W19865, W17012);
not G21563 (W20166, W20168);
or G21564 (W20167, W20290, W17714);
not G21565 (W20168, W20291);
and G21566 (W20169, W19864, W17682);
not G21567 (W20170, W14569);
and G21568 (W20171, W12911, W18961);
and G21569 (W20172, W17682, W15630, W18961);
not G21570 (W20173, W14569);
nand G21571 (W20174, W16982, W10575);
nand G21572 (W20175, W16950, W20292);
nand G21573 (W20176, W10563, W20292);
nand G21574 (W20177, W16994, W20293);
nand G21575 (W20178, W10587, W20293);
nand G21576 (W20179, W17000, W10555);
nand G21577 (W20180, W16957, W10571);
nand G21578 (W20181, W16964, W10583);
nand G21579 (W20182, W16978, W20294);
nand G21580 (W20183, W10567, W20294);
nand G21581 (W20184, W16968, W20295);
nand G21582 (W20185, W10551, W20295);
nand G21583 (W20186, W16974, W10559);
nand G21584 (W20187, W16986, W10579);
or G21585 (W20188, W19452, W19877, W19455);
or G21586 (W20189, W19461, W19885, W19464);
not G21587 (W20190, W20191);
not G21588 (W20191, W20296);
not G21589 (W20192, W20193);
not G21590 (W20193, W20297);
not G21591 (W20194, W20195);
not G21592 (W20195, W20298);
not G21593 (W20196, W20197);
not G21594 (W20197, W20299);
not G21595 (W20198, W17795);
not G21596 (W20199, W17795);
not G21597 (W20200, W17795);
not G21598 (W20201, W17795);
not G21599 (W20202, W17795);
nand G21600 (W20203, W19943, W19944, W17167);
not G21601 (W20204, W20206);
or G21602 (W20205, W20300, W17861);
not G21603 (W20206, W20301);
and G21604 (W20207, W19943, W17829);
not G21605 (W20208, W14840);
and G21606 (W20209, W13306, W19063);
and G21607 (W20210, W17829, W15812, W19063);
not G21608 (W20211, W14840);
nand G21609 (W20212, W17137, W11344);
nand G21610 (W20213, W17105, W20302);
nand G21611 (W20214, W11332, W20302);
nand G21612 (W20215, W17149, W20303);
nand G21613 (W20216, W11356, W20303);
nand G21614 (W20217, W17155, W11324);
nand G21615 (W20218, W17112, W11340);
nand G21616 (W20219, W17119, W11352);
nand G21617 (W20220, W17133, W20304);
nand G21618 (W20221, W11336, W20304);
nand G21619 (W20222, W17123, W20305);
nand G21620 (W20223, W11363, W20305);
nand G21621 (W20224, W17129, W11328);
nand G21622 (W20225, W17141, W11348);
or G21623 (W20226, W19543, W19956, W19546);
or G21624 (W20227, W19552, W19964, W19555);
not G21625 (W20228, W20306);
not G21626 (W20229, W8613);
not G21627 (W20230, W8616);
not G21628 (W20231, W9386);
not G21629 (W20232, W9389);
not G21630 (W20233, W8609);
not G21631 (W20234, W10159);
not G21632 (W20235, W10162);
not G21633 (W20236, W9382);
nand G21634 (W20237, W20239, W20249);
nand G21635 (W20238, W20307, W20249);
nor G21636 (W20239, W19994, W20264, W20308, W20309);
not G21637 (W20240, I1633);
not G21638 (W20241, I1634);
not G21639 (W20242, I1635);
not G21640 (W20243, I1636);
not G21641 (W20244, I1637);
not G21642 (W20245, I1638);
not G21643 (W20246, W20310);
not G21644 (W20247, W20311);
nor G21645 (W20248, W20265, W20264, W19996, W20309);
not G21646 (W20249, W20312);
nor G21647 (W20250, W19994, W19995, W19996, W20309);
nor G21648 (W20251, W20265, W19995, W19996, W20309);
nor G21649 (W20252, W19994, W20264, W20308, W19997);
nor G21650 (W20253, W19994, W19995, W20308, W19997);
nor G21651 (W20254, W19994, W20264, W19996, W20309);
not G21652 (W20255, W20313);
nand G21653 (W20256, W19592, W20249);
nand G21654 (W20257, W20314, W20249);
nand G21655 (W20258, W20026, W20249);
nand G21656 (W20259, W20027, W20249);
nand G21657 (W20260, W20315, W20249);
nand G21658 (W20261, W20316, W20249);
not G21659 (W20262, W20317);
nor G21660 (W20263, W20265, W20264, W20308, W19997);
not G21661 (W20264, W20318);
not G21662 (W20265, I1633);
not G21663 (W20266, W17356);
not G21664 (W20267, W17356);
not G21665 (W20268, W17356);
not G21666 (W20269, W17356);
not G21667 (W20270, W20319);
not G21668 (W20271, W13982);
nand G21669 (W20272, W16640, W9021);
nand G21670 (W20273, W16684, W9005);
nand G21671 (W20274, W16668, W9025);
nand G21672 (W20275, W16658, W9009);
not G21673 (W20276, W17502);
not G21674 (W20277, W17502);
not G21675 (W20278, W17502);
not G21676 (W20279, W17502);
not G21677 (W20280, W20320);
not G21678 (W20281, W14276);
nand G21679 (W20282, W16795, W9794);
nand G21680 (W20283, W16839, W9778);
nand G21681 (W20284, W16823, W9798);
nand G21682 (W20285, W16813, W9782);
not G21683 (W20286, W17648);
not G21684 (W20287, W17648);
not G21685 (W20288, W17648);
not G21686 (W20289, W17648);
not G21687 (W20290, W20321);
not G21688 (W20291, W14569);
nand G21689 (W20292, W16950, W10563);
nand G21690 (W20293, W16994, W10587);
nand G21691 (W20294, W16978, W10567);
nand G21692 (W20295, W16968, W10551);
not G21693 (W20296, W17795);
not G21694 (W20297, W17795);
not G21695 (W20298, W17795);
not G21696 (W20299, W17795);
not G21697 (W20300, W20322);
not G21698 (W20301, W14840);
nand G21699 (W20302, W17105, W11332);
nand G21700 (W20303, W17149, W11356);
nand G21701 (W20304, W17133, W11336);
nand G21702 (W20305, W17123, W11363);
not G21703 (W20306, W20323);
nor G21704 (W20307, W20265, W19995, W19996, W19997);
not G21705 (W20308, I1634);
not G21706 (W20309, W20324);
not G21707 (W20310, I1639);
not G21708 (W20311, W20325);
not G21709 (W20312, W20326);
nor G21710 (W20313, I1640, I1641);
nor G21711 (W20314, W20265, W19995, W20308, W20309);
nor G21712 (W20315, W20265, W20264, W20308, W20309);
nor G21713 (W20316, W19994, W19995, W20308, W20309);
nand G21714 (W20317, W20327, W20328);
not G21715 (W20318, I1579);
nand G21716 (W20319, W15194, W19288, W9108);
nand G21717 (W20320, W15388, W19379, W9881);
nand G21718 (W20321, W15581, W19470, W10654);
nand G21719 (W20322, W15763, W19561, W11427);
nor G21720 (W20323, I1642, I1643);
not G21721 (W20324, I1580);
not G21722 (W20325, I1644);
nor G21723 (W20326, I1635, W20243, I1637, I1638);
or G21724 (W20327, W20329, W20008);
or G21725 (W20328, W20330, W20228);
not G21726 (W20329, I1568);
not G21727 (W20330, I1571);
endmodule