
module aes_sbox ( a, d );
  input [7:0] a;
  output [7:0] d;
  wire   n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626,
         n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636,
         n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646,
         n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656,
         n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666,
         n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676,
         n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686,
         n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696,
         n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706,
         n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716,
         n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726,
         n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736,
         n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746,
         n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756,
         n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766,
         n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776,
         n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786,
         n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796,
         n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806,
         n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816,
         n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826,
         n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836,
         n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846,
         n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856,
         n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866,
         n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876,
         n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886,
         n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896,
         n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906,
         n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916,
         n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926,
         n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936,
         n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946,
         n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956,
         n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966,
         n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976,
         n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986,
         n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996,
         n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006,
         n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016,
         n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026,
         n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036,
         n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046,
         n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056,
         n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066,
         n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076,
         n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086,
         n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096,
         n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106,
         n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116,
         n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126,
         n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136,
         n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146,
         n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156,
         n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166,
         n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176,
         n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186,
         n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196,
         n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206,
         n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216,
         n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226,
         n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236,
         n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246,
         n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256,
         n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266,
         n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276,
         n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286,
         n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296,
         n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306,
         n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316,
         n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326,
         n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336,
         n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346,
         n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356,
         n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366,
         n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376,
         n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386,
         n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396,
         n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406,
         n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416,
         n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426,
         n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436,
         n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446,
         n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456,
         n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466,
         n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476,
         n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486,
         n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496,
         n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506,
         n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516,
         n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526,
         n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536,
         n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546,
         n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556,
         n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566,
         n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576,
         n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586,
         n3587, n3588;

  OR2X1TS U1658 ( .A(n3556), .B(n3563), .Y(n3202) );
  NOR2X1TS U1659 ( .A(n2716), .B(n2819), .Y(n2617) );
  NAND2X1TS U1660 ( .A(n2851), .B(n2744), .Y(n2618) );
  NAND2X1TS U1661 ( .A(n3391), .B(n2618), .Y(n2619) );
  NOR2X1TS U1662 ( .A(n2617), .B(n2619), .Y(n2620) );
  NAND2X1TS U1663 ( .A(n3018), .B(n2620), .Y(n2621) );
  NOR2X1TS U1664 ( .A(n2838), .B(n2774), .Y(n2622) );
  NOR2X1TS U1665 ( .A(n2771), .B(n2768), .Y(n2623) );
  NOR2X1TS U1666 ( .A(n3222), .B(n2704), .Y(n2624) );
  NOR2X1TS U1667 ( .A(n2782), .B(n2815), .Y(n2625) );
  NOR2X1TS U1668 ( .A(n2622), .B(n2623), .Y(n2626) );
  NOR2X1TS U1669 ( .A(n2624), .B(n2625), .Y(n2627) );
  NAND2X1TS U1670 ( .A(n2626), .B(n2627), .Y(n2628) );
  NOR2X1TS U1671 ( .A(n3357), .B(n3358), .Y(n2629) );
  NAND2X1TS U1672 ( .A(n3085), .B(n3356), .Y(n2630) );
  NAND2X1TS U1673 ( .A(n2629), .B(n2630), .Y(n2631) );
  NOR2X1TS U1674 ( .A(n2628), .B(n2631), .Y(n2632) );
  NAND2X1TS U1675 ( .A(n3017), .B(n2632), .Y(n2633) );
  NOR2X1TS U1676 ( .A(n2621), .B(n2633), .Y(n2634) );
  NAND2X1TS U1677 ( .A(n2965), .B(n2634), .Y(n2635) );
  NOR2BX1TS U1678 ( .AN(n2955), .B(n2635), .Y(n3060) );
  NAND2X1TS U1679 ( .A(n2877), .B(n2784), .Y(n2636) );
  NAND2X1TS U1680 ( .A(n3391), .B(n2636), .Y(n2637) );
  NOR2X1TS U1681 ( .A(n3462), .B(n3463), .Y(n2638) );
  NOR2X1TS U1682 ( .A(n2894), .B(n3461), .Y(n2639) );
  NAND2X1TS U1683 ( .A(n2871), .B(n2639), .Y(n2640) );
  NAND2X1TS U1684 ( .A(n2638), .B(n2640), .Y(n2641) );
  NAND2X1TS U1685 ( .A(n3004), .B(n3458), .Y(n2642) );
  NAND2X1TS U1686 ( .A(n3114), .B(n2642), .Y(n2643) );
  NOR2X1TS U1687 ( .A(n2831), .B(n2982), .Y(n2644) );
  NOR2X1TS U1688 ( .A(n2788), .B(n2990), .Y(n2645) );
  NOR2X1TS U1689 ( .A(n2641), .B(n2643), .Y(n2646) );
  NOR2X1TS U1690 ( .A(n2644), .B(n2645), .Y(n2647) );
  NAND2X1TS U1691 ( .A(n2646), .B(n2647), .Y(n2648) );
  NOR2X1TS U1692 ( .A(n2794), .B(n3095), .Y(n2649) );
  NOR2X1TS U1693 ( .A(n2637), .B(n2648), .Y(n2650) );
  NOR2X1TS U1694 ( .A(n3176), .B(n2649), .Y(n2651) );
  NAND2X1TS U1695 ( .A(n2650), .B(n2651), .Y(n2652) );
  NAND2BX1TS U1696 ( .AN(n2652), .B(n3248), .Y(n2653) );
  NOR2X1TS U1697 ( .A(n3053), .B(n2653), .Y(n2654) );
  NAND2X1TS U1698 ( .A(n3164), .B(n2654), .Y(d[0]) );
  AND2X1TS U1699 ( .A(n3428), .B(n3500), .Y(n3141) );
  NOR2BX1TS U1700 ( .AN(n3248), .B(n3165), .Y(n2655) );
  NAND2X1TS U1701 ( .A(n2787), .B(n2778), .Y(n2656) );
  NAND2X1TS U1702 ( .A(n3115), .B(n2737), .Y(n2657) );
  NAND2X1TS U1703 ( .A(n2656), .B(n2657), .Y(n2658) );
  NAND2X1TS U1704 ( .A(n3220), .B(n3219), .Y(n2659) );
  NOR2X1TS U1705 ( .A(n3223), .B(n3224), .Y(n2660) );
  NAND2X1TS U1706 ( .A(n2745), .B(n3221), .Y(n2661) );
  NAND2X1TS U1707 ( .A(n2660), .B(n2661), .Y(n2662) );
  NOR2X1TS U1708 ( .A(n2833), .B(n2807), .Y(n2663) );
  AND2X1TS U1709 ( .A(n2846), .B(n2748), .Y(n2664) );
  NOR2X1TS U1710 ( .A(n2659), .B(n2662), .Y(n2665) );
  NOR2X1TS U1711 ( .A(n2663), .B(n2664), .Y(n2666) );
  NAND2X1TS U1712 ( .A(n2665), .B(n2666), .Y(n2667) );
  NOR2X1TS U1713 ( .A(n2658), .B(n2667), .Y(n2668) );
  NAND2X1TS U1714 ( .A(n3031), .B(n2668), .Y(n2669) );
  NOR2X1TS U1715 ( .A(n2669), .B(n3179), .Y(n2670) );
  NOR2X1TS U1716 ( .A(n3196), .B(n3203), .Y(n2671) );
  NAND2X1TS U1717 ( .A(n2670), .B(n2671), .Y(n2672) );
  NOR2X1TS U1718 ( .A(n3247), .B(n2672), .Y(n2673) );
  NAND2X1TS U1719 ( .A(n2655), .B(n2673), .Y(d[2]) );
  NOR2X1TS U1720 ( .A(n2840), .B(n3171), .Y(n2674) );
  NOR2X1TS U1721 ( .A(n2830), .B(n2712), .Y(n2675) );
  NOR2X1TS U1722 ( .A(n2674), .B(n2675), .Y(n2676) );
  NAND2X1TS U1723 ( .A(n2851), .B(n2779), .Y(n2677) );
  NAND2X1TS U1724 ( .A(n2676), .B(n2677), .Y(n2678) );
  NAND2X1TS U1725 ( .A(n2726), .B(n3170), .Y(n2679) );
  NAND2X1TS U1726 ( .A(n2785), .B(n3166), .Y(n2680) );
  NAND2X1TS U1727 ( .A(n2679), .B(n2680), .Y(n2681) );
  NOR2BX1TS U1728 ( .AN(n2849), .B(n3167), .Y(n2682) );
  NOR2X1TS U1729 ( .A(n2682), .B(n2681), .Y(n2683) );
  NAND2X1TS U1730 ( .A(n2933), .B(n3168), .Y(n2684) );
  NAND2X1TS U1731 ( .A(n2683), .B(n2684), .Y(n2685) );
  NOR2X1TS U1732 ( .A(n2719), .B(n2761), .Y(n2686) );
  NOR2X1TS U1733 ( .A(n3172), .B(n2686), .Y(n2687) );
  NAND2X1TS U1734 ( .A(n3070), .B(n2687), .Y(n2688) );
  NOR2X1TS U1735 ( .A(n2678), .B(n2685), .Y(n2689) );
  NOR2X1TS U1736 ( .A(n2688), .B(n3165), .Y(n2690) );
  NAND2X1TS U1737 ( .A(n2689), .B(n2690), .Y(n2691) );
  NOR2X1TS U1738 ( .A(n3028), .B(n2691), .Y(n2692) );
  NAND2X1TS U1739 ( .A(n3164), .B(n2692), .Y(d[3]) );
  AND2X2TS U1740 ( .A(n3500), .B(n3555), .Y(n2693) );
  AND2X2TS U1741 ( .A(n2706), .B(n3555), .Y(n2694) );
  AND2X2TS U1742 ( .A(n3500), .B(n3460), .Y(n2695) );
  AND2X2TS U1743 ( .A(n2913), .B(n3446), .Y(n2696) );
  OR2X2TS U1744 ( .A(n3568), .B(n3569), .Y(n2697) );
  AND2X2TS U1745 ( .A(n3446), .B(n3562), .Y(n2698) );
  AND2X2TS U1746 ( .A(n2903), .B(n3304), .Y(n2699) );
  AND2X2TS U1747 ( .A(n3499), .B(n3459), .Y(n2700) );
  AND2X2TS U1748 ( .A(n3370), .B(n3466), .Y(n2701) );
  OR2X2TS U1749 ( .A(n2863), .B(n2857), .Y(n2702) );
  NAND2X1TS U1750 ( .A(n2905), .B(n2893), .Y(n2703) );
  INVXLTS U1751 ( .A(n2994), .Y(n2704) );
  INVXLTS U1752 ( .A(n2994), .Y(n2705) );
  INVXLTS U1753 ( .A(n2703), .Y(n2706) );
  INVXLTS U1754 ( .A(n2703), .Y(n2707) );
  INVXLTS U1755 ( .A(n3460), .Y(n2708) );
  INVXLTS U1756 ( .A(n2708), .Y(n2709) );
  INVXLTS U1757 ( .A(n2933), .Y(n2710) );
  INVXLTS U1758 ( .A(n2702), .Y(n2711) );
  INVXLTS U1759 ( .A(n2702), .Y(n2712) );
  INVXLTS U1760 ( .A(n3096), .Y(n2713) );
  INVXLTS U1761 ( .A(n3096), .Y(n2714) );
  INVXLTS U1762 ( .A(n2939), .Y(n2715) );
  INVXLTS U1763 ( .A(n2939), .Y(n2716) );
  INVXLTS U1764 ( .A(n3131), .Y(n2717) );
  INVXLTS U1765 ( .A(n3131), .Y(n2718) );
  INVXLTS U1766 ( .A(n2925), .Y(n2719) );
  INVXLTS U1767 ( .A(n2925), .Y(n2720) );
  INVXLTS U1768 ( .A(n2975), .Y(n2721) );
  INVXLTS U1769 ( .A(n2975), .Y(n2722) );
  INVXLTS U1770 ( .A(n2700), .Y(n2723) );
  INVXLTS U1771 ( .A(n2700), .Y(n2724) );
  INVXLTS U1772 ( .A(n3202), .Y(n2725) );
  INVXLTS U1773 ( .A(n3202), .Y(n2726) );
  INVXLTS U1774 ( .A(n2935), .Y(n2727) );
  INVXLTS U1775 ( .A(n2935), .Y(n2728) );
  INVXLTS U1776 ( .A(n2697), .Y(n2729) );
  INVXLTS U1777 ( .A(n2697), .Y(n2730) );
  INVXLTS U1778 ( .A(n2699), .Y(n2731) );
  INVXLTS U1779 ( .A(n2699), .Y(n2732) );
  INVXLTS U1780 ( .A(n2698), .Y(n2733) );
  INVXLTS U1781 ( .A(n2698), .Y(n2734) );
  INVXLTS U1782 ( .A(n3161), .Y(n2735) );
  INVXLTS U1783 ( .A(n3161), .Y(n2736) );
  INVXLTS U1784 ( .A(n3080), .Y(n2737) );
  INVXLTS U1785 ( .A(n3080), .Y(n2738) );
  INVXLTS U1786 ( .A(n2701), .Y(n2739) );
  INVXLTS U1787 ( .A(n2701), .Y(n2740) );
  INVXLTS U1788 ( .A(n2945), .Y(n2741) );
  INVXLTS U1789 ( .A(n2741), .Y(n2742) );
  INVXLTS U1790 ( .A(n2741), .Y(n2743) );
  INVXLTS U1791 ( .A(n2945), .Y(n2744) );
  INVXLTS U1792 ( .A(n2945), .Y(n2745) );
  INVXLTS U1793 ( .A(n3006), .Y(n2746) );
  INVXLTS U1794 ( .A(n2746), .Y(n2747) );
  INVXLTS U1795 ( .A(n2746), .Y(n2748) );
  INVXLTS U1796 ( .A(n3023), .Y(n2749) );
  INVXLTS U1797 ( .A(n2749), .Y(n2750) );
  INVXLTS U1798 ( .A(n2988), .Y(n2751) );
  INVXLTS U1799 ( .A(n2751), .Y(n2752) );
  INVXLTS U1800 ( .A(n2751), .Y(n2753) );
  INVXLTS U1801 ( .A(n3089), .Y(n2754) );
  INVXLTS U1802 ( .A(n3089), .Y(n2756) );
  INVXLTS U1803 ( .A(n3089), .Y(n2755) );
  INVXLTS U1804 ( .A(n2928), .Y(n2757) );
  INVXLTS U1805 ( .A(n2928), .Y(n2759) );
  INVXLTS U1806 ( .A(n2928), .Y(n2758) );
  INVXLTS U1807 ( .A(n2693), .Y(n2760) );
  INVXLTS U1808 ( .A(n2693), .Y(n2762) );
  INVXLTS U1809 ( .A(n2693), .Y(n2761) );
  INVXLTS U1810 ( .A(n3125), .Y(n2763) );
  INVXLTS U1811 ( .A(n3125), .Y(n2765) );
  INVXLTS U1812 ( .A(n3125), .Y(n2764) );
  INVXLTS U1813 ( .A(n2986), .Y(n2766) );
  INVXLTS U1814 ( .A(n2986), .Y(n2768) );
  INVXLTS U1815 ( .A(n2986), .Y(n2767) );
  INVXLTS U1816 ( .A(n2760), .Y(n2769) );
  INVXLTS U1817 ( .A(n2762), .Y(n2770) );
  INVXLTS U1818 ( .A(n3051), .Y(n2772) );
  INVXLTS U1819 ( .A(n3051), .Y(n2771) );
  INVXLTS U1820 ( .A(n3013), .Y(n2773) );
  INVXLTS U1821 ( .A(n2773), .Y(n2774) );
  INVXLTS U1822 ( .A(n2773), .Y(n2776) );
  INVXLTS U1823 ( .A(n2773), .Y(n2775) );
  INVXLTS U1824 ( .A(n3085), .Y(n2777) );
  INVXLTS U1825 ( .A(n2777), .Y(n2778) );
  INVXLTS U1826 ( .A(n2777), .Y(n2779) );
  INVXLTS U1827 ( .A(n3077), .Y(n2780) );
  INVXLTS U1828 ( .A(n3077), .Y(n2782) );
  INVXLTS U1829 ( .A(n3077), .Y(n2781) );
  INVXLTS U1830 ( .A(n2791), .Y(n2783) );
  INVXLTS U1831 ( .A(n2793), .Y(n2784) );
  INVXLTS U1832 ( .A(n3013), .Y(n2785) );
  INVXLTS U1833 ( .A(n3013), .Y(n2787) );
  INVXLTS U1834 ( .A(n3013), .Y(n2786) );
  INVXLTS U1835 ( .A(n2763), .Y(n2788) );
  INVXLTS U1836 ( .A(n2765), .Y(n2790) );
  INVXLTS U1837 ( .A(n2764), .Y(n2789) );
  INVXLTS U1838 ( .A(n2695), .Y(n2791) );
  INVXLTS U1839 ( .A(n2695), .Y(n2793) );
  INVXLTS U1840 ( .A(n2695), .Y(n2792) );
  INVXLTS U1841 ( .A(n2694), .Y(n2794) );
  INVXLTS U1842 ( .A(n2694), .Y(n2796) );
  INVXLTS U1843 ( .A(n2694), .Y(n2795) );
  INVXLTS U1844 ( .A(n2988), .Y(n2798) );
  INVXLTS U1845 ( .A(n2988), .Y(n2797) );
  INVXLTS U1846 ( .A(n3015), .Y(n2799) );
  INVXLTS U1847 ( .A(n2799), .Y(n2800) );
  INVXLTS U1848 ( .A(n2799), .Y(n2801) );
  INVXLTS U1849 ( .A(n3141), .Y(n2802) );
  INVXLTS U1850 ( .A(n3141), .Y(n2804) );
  INVXLTS U1851 ( .A(n3141), .Y(n2803) );
  INVXLTS U1852 ( .A(n2946), .Y(n2805) );
  INVXLTS U1853 ( .A(n2946), .Y(n2807) );
  INVXLTS U1854 ( .A(n2946), .Y(n2806) );
  INVXLTS U1855 ( .A(n2699), .Y(n2808) );
  INVXLTS U1856 ( .A(n2808), .Y(n2809) );
  INVXLTS U1857 ( .A(n2808), .Y(n2811) );
  INVXLTS U1858 ( .A(n2808), .Y(n2810) );
  INVXLTS U1859 ( .A(n3096), .Y(n2812) );
  INVXLTS U1860 ( .A(n2812), .Y(n2813) );
  INVXLTS U1861 ( .A(n2812), .Y(n2815) );
  INVXLTS U1862 ( .A(n2812), .Y(n2814) );
  INVXLTS U1863 ( .A(n2796), .Y(n2816) );
  INVXLTS U1864 ( .A(n2794), .Y(n2817) );
  INVXLTS U1865 ( .A(n3131), .Y(n2818) );
  INVXLTS U1866 ( .A(n2818), .Y(n2819) );
  INVXLTS U1867 ( .A(n2818), .Y(n2821) );
  INVXLTS U1868 ( .A(n2818), .Y(n2820) );
  INVXLTS U1869 ( .A(n2696), .Y(n2822) );
  INVXLTS U1870 ( .A(n2696), .Y(n2824) );
  INVXLTS U1871 ( .A(n2696), .Y(n2823) );
  INVXLTS U1872 ( .A(n3080), .Y(n2825) );
  INVXLTS U1873 ( .A(n2825), .Y(n2826) );
  INVXLTS U1874 ( .A(n2825), .Y(n2828) );
  INVXLTS U1875 ( .A(n2825), .Y(n2827) );
  INVXLTS U1876 ( .A(n2755), .Y(n2829) );
  INVXLTS U1877 ( .A(n2756), .Y(n2830) );
  INVXLTS U1878 ( .A(n2754), .Y(n2831) );
  INVXLTS U1879 ( .A(n3202), .Y(n2832) );
  INVXLTS U1880 ( .A(n2832), .Y(n2835) );
  INVXLTS U1881 ( .A(n2832), .Y(n2833) );
  INVXLTS U1882 ( .A(n2832), .Y(n2834) );
  INVXLTS U1883 ( .A(n2954), .Y(n2836) );
  INVXLTS U1884 ( .A(n2836), .Y(n2837) );
  INVXLTS U1885 ( .A(n2836), .Y(n2838) );
  INVXLTS U1886 ( .A(n2836), .Y(n2839) );
  INVXLTS U1887 ( .A(n3051), .Y(n2840) );
  INVXLTS U1888 ( .A(n2840), .Y(n2841) );
  INVXLTS U1889 ( .A(n2840), .Y(n2842) );
  INVXLTS U1890 ( .A(n2700), .Y(n2843) );
  INVXLTS U1891 ( .A(n2843), .Y(n2844) );
  INVXLTS U1892 ( .A(n2843), .Y(n2846) );
  INVXLTS U1893 ( .A(n2843), .Y(n2845) );
  INVXLTS U1894 ( .A(n2946), .Y(n2847) );
  INVXLTS U1895 ( .A(n2847), .Y(n2848) );
  INVXLTS U1896 ( .A(n2847), .Y(n2849) );
  INVXLTS U1897 ( .A(n3141), .Y(n2850) );
  INVXLTS U1898 ( .A(n2850), .Y(n2851) );
  INVXLTS U1899 ( .A(n2850), .Y(n2852) );
  INVXLTS U1900 ( .A(n3161), .Y(n2853) );
  INVXLTS U1901 ( .A(n2853), .Y(n2854) );
  INVXLTS U1902 ( .A(n2853), .Y(n2855) );
  INVXLTS U1903 ( .A(n2939), .Y(n2856) );
  INVXLTS U1904 ( .A(n2856), .Y(n2857) );
  INVXLTS U1905 ( .A(n2856), .Y(n2858) );
  INVXLTS U1906 ( .A(n2767), .Y(n2859) );
  INVXLTS U1907 ( .A(n2766), .Y(n2860) );
  INVXLTS U1908 ( .A(n2933), .Y(n2861) );
  INVXLTS U1909 ( .A(n2861), .Y(n2862) );
  INVXLTS U1910 ( .A(n2861), .Y(n2863) );
  INVXLTS U1911 ( .A(n3077), .Y(n2864) );
  INVXLTS U1912 ( .A(n2864), .Y(n2865) );
  INVXLTS U1913 ( .A(n2864), .Y(n2867) );
  INVXLTS U1914 ( .A(n2864), .Y(n2866) );
  INVXLTS U1915 ( .A(n2975), .Y(n2868) );
  INVXLTS U1916 ( .A(n2868), .Y(n2869) );
  INVXLTS U1917 ( .A(n2868), .Y(n2871) );
  INVXLTS U1918 ( .A(n2868), .Y(n2870) );
  INVXLTS U1919 ( .A(n2994), .Y(n2872) );
  INVXLTS U1920 ( .A(n2872), .Y(n2873) );
  INVXLTS U1921 ( .A(n2872), .Y(n2874) );
  INVXLTS U1922 ( .A(n2872), .Y(n2875) );
  INVXLTS U1923 ( .A(n2928), .Y(n2876) );
  INVXLTS U1924 ( .A(n2876), .Y(n2877) );
  INVXLTS U1925 ( .A(n2876), .Y(n2878) );
  INVXLTS U1926 ( .A(n2876), .Y(n2879) );
  INVXLTS U1927 ( .A(n2925), .Y(n2880) );
  INVXLTS U1928 ( .A(n2880), .Y(n2881) );
  INVXLTS U1929 ( .A(n2880), .Y(n2882) );
  INVXLTS U1930 ( .A(n2880), .Y(n2883) );
  INVXLTS U1931 ( .A(n2935), .Y(n2884) );
  INVXLTS U1932 ( .A(n2884), .Y(n2885) );
  INVXLTS U1933 ( .A(n2884), .Y(n2888) );
  INVXLTS U1934 ( .A(n2884), .Y(n2886) );
  INVXLTS U1935 ( .A(n2884), .Y(n2887) );
  INVXLTS U1936 ( .A(a[2]), .Y(n2889) );
  INVXLTS U1937 ( .A(n2889), .Y(n2890) );
  INVXLTS U1938 ( .A(n2889), .Y(n2891) );
  INVXLTS U1939 ( .A(a[7]), .Y(n2892) );
  INVXLTS U1940 ( .A(n2892), .Y(n2893) );
  INVXLTS U1941 ( .A(n2892), .Y(n2894) );
  INVXLTS U1942 ( .A(a[6]), .Y(n2895) );
  INVXLTS U1943 ( .A(n2895), .Y(n2896) );
  INVXLTS U1944 ( .A(n2895), .Y(n2897) );
  INVXLTS U1945 ( .A(a[3]), .Y(n2898) );
  INVXLTS U1946 ( .A(n2898), .Y(n2899) );
  INVXLTS U1947 ( .A(n2898), .Y(n2900) );
  INVXLTS U1948 ( .A(a[0]), .Y(n2901) );
  INVXLTS U1949 ( .A(n2901), .Y(n2902) );
  INVXLTS U1950 ( .A(n2901), .Y(n2903) );
  INVXLTS U1951 ( .A(a[5]), .Y(n2904) );
  INVXLTS U1952 ( .A(n2904), .Y(n2905) );
  INVXLTS U1953 ( .A(n2904), .Y(n2906) );
  INVXLTS U1954 ( .A(a[4]), .Y(n2907) );
  INVXLTS U1955 ( .A(n2907), .Y(n2908) );
  INVXLTS U1956 ( .A(n2907), .Y(n2909) );
  INVXLTS U1957 ( .A(a[1]), .Y(n2910) );
  INVXLTS U1958 ( .A(n2910), .Y(n2911) );
  INVXLTS U1959 ( .A(n2910), .Y(n2913) );
  INVXLTS U1960 ( .A(n2910), .Y(n2912) );
  AND2XLTS U1961 ( .A(n2718), .B(n3464), .Y(n3463) );
  NOR2XLTS U1962 ( .A(n2736), .B(n3465), .Y(n3462) );
  NOR2XLTS U1963 ( .A(n2963), .B(n2964), .Y(n2962) );
  NOR2XLTS U1964 ( .A(n2967), .B(n2968), .Y(n2966) );
  NOR2XLTS U1965 ( .A(n2971), .B(n2972), .Y(n2970) );
  NOR2XLTS U1966 ( .A(n2977), .B(n2734), .Y(n2971) );
  NOR2XLTS U1967 ( .A(n2978), .B(n2979), .Y(n2969) );
  NOR2XLTS U1968 ( .A(n2750), .B(n2745), .Y(n2990) );
  NOR2XLTS U1969 ( .A(n2917), .B(n2991), .Y(n2961) );
  NOR2XLTS U1970 ( .A(n3028), .B(n3029), .Y(n3027) );
  NOR2XLTS U1971 ( .A(n3032), .B(n3033), .Y(n3030) );
  NOR2XLTS U1972 ( .A(n3036), .B(n3037), .Y(n3035) );
  NOR2XLTS U1973 ( .A(n2734), .B(n2772), .Y(n3037) );
  NOR2XLTS U1974 ( .A(n3038), .B(n3039), .Y(n3034) );
  NOR2XLTS U1975 ( .A(n2711), .B(n2735), .Y(n3039) );
  NOR2XLTS U1976 ( .A(n3040), .B(n2805), .Y(n3038) );
  NOR2XLTS U1977 ( .A(n3043), .B(n3044), .Y(n3042) );
  AND2XLTS U1978 ( .A(n2846), .B(n2976), .Y(n3044) );
  NOR2XLTS U1979 ( .A(n2891), .B(n2913), .Y(n3046) );
  NOR2XLTS U1980 ( .A(n3047), .B(n2710), .Y(n3043) );
  NOR2XLTS U1981 ( .A(n3048), .B(n3049), .Y(n3041) );
  NOR2XLTS U1982 ( .A(n3050), .B(n2739), .Y(n3049) );
  NOR2XLTS U1983 ( .A(n2694), .B(n2841), .Y(n3050) );
  NOR2XLTS U1984 ( .A(n2839), .B(n2947), .Y(n3048) );
  NOR2XLTS U1985 ( .A(n3052), .B(n3053), .Y(n3026) );
  OR2XLTS U1986 ( .A(n3203), .B(n3467), .Y(n3053) );
  NOR2XLTS U1987 ( .A(n3470), .B(n3471), .Y(n3469) );
  NOR2XLTS U1988 ( .A(n2831), .B(n2824), .Y(n3470) );
  NOR2XLTS U1989 ( .A(n3474), .B(n3475), .Y(n3468) );
  NOR2XLTS U1990 ( .A(n3483), .B(n3484), .Y(n3479) );
  NOR2XLTS U1991 ( .A(n3485), .B(n2821), .Y(n3484) );
  NOR2XLTS U1992 ( .A(n2858), .B(n2878), .Y(n3485) );
  NOR2XLTS U1993 ( .A(n3486), .B(n2760), .Y(n3483) );
  NOR2XLTS U1994 ( .A(n2867), .B(n3446), .Y(n3486) );
  NOR2XLTS U1995 ( .A(n3056), .B(n3057), .Y(n3055) );
  NOR2XLTS U1996 ( .A(n2804), .B(n2758), .Y(n3056) );
  NOR2XLTS U1997 ( .A(n3058), .B(n3059), .Y(n3054) );
  NOR2XLTS U1998 ( .A(n2963), .B(n3062), .Y(n3061) );
  NOR2XLTS U1999 ( .A(n3067), .B(n3068), .Y(n3066) );
  NOR2XLTS U2000 ( .A(n2837), .B(n2806), .Y(n3067) );
  NOR2XLTS U2001 ( .A(n3098), .B(n3099), .Y(n3063) );
  NOR2XLTS U2002 ( .A(n3107), .B(n3108), .Y(n3106) );
  NOR2XLTS U2003 ( .A(n3109), .B(n2781), .Y(n3108) );
  NOR2XLTS U2004 ( .A(n3110), .B(n2804), .Y(n3107) );
  NOR2XLTS U2005 ( .A(n3111), .B(n3112), .Y(n3105) );
  NOR2XLTS U2006 ( .A(n2719), .B(n2732), .Y(n3111) );
  OR2XLTS U2007 ( .A(n2953), .B(n3116), .Y(n2963) );
  NOR2XLTS U2008 ( .A(n3119), .B(n3120), .Y(n3118) );
  NOR2XLTS U2009 ( .A(n3123), .B(n3124), .Y(n3122) );
  NOR2XLTS U2010 ( .A(n2705), .B(n2790), .Y(n3124) );
  NOR2XLTS U2011 ( .A(n3126), .B(n3127), .Y(n3121) );
  NOR2XLTS U2012 ( .A(n3133), .B(n2735), .Y(n3126) );
  NOR2XLTS U2013 ( .A(n2888), .B(n3134), .Y(n3133) );
  NOR2XLTS U2014 ( .A(n3135), .B(n2815), .Y(n3119) );
  NOR2XLTS U2015 ( .A(n3023), .B(n3136), .Y(n3135) );
  NOR2XLTS U2016 ( .A(n3137), .B(n3138), .Y(n3117) );
  NOR2XLTS U2017 ( .A(n2916), .B(n2917), .Y(n2915) );
  NOR2XLTS U2018 ( .A(n2997), .B(n2998), .Y(n2996) );
  NOR2XLTS U2019 ( .A(n3001), .B(n3002), .Y(n3000) );
  NOR2XLTS U2020 ( .A(n2977), .B(n3003), .Y(n3002) );
  NOR2XLTS U2021 ( .A(n3005), .B(n2736), .Y(n3001) );
  NOR2XLTS U2022 ( .A(n2881), .B(n2748), .Y(n3005) );
  NOR2XLTS U2023 ( .A(n3007), .B(n3008), .Y(n2999) );
  NOR2XLTS U2024 ( .A(n3011), .B(n3012), .Y(n3009) );
  NOR2XLTS U2025 ( .A(n2776), .B(n2743), .Y(n3012) );
  NOR2XLTS U2026 ( .A(n3014), .B(n2801), .Y(n3011) );
  NOR2XLTS U2027 ( .A(n3016), .B(n2822), .Y(n3007) );
  NOR2XLTS U2028 ( .A(n3019), .B(n3020), .Y(n2995) );
  NOR2XLTS U2029 ( .A(n3024), .B(n3025), .Y(n3021) );
  NOR2XLTS U2030 ( .A(n2759), .B(n2771), .Y(n3025) );
  NOR2XLTS U2031 ( .A(n2954), .B(n2724), .Y(n3024) );
  NOR2XLTS U2032 ( .A(n2920), .B(n2921), .Y(n2919) );
  NOR2XLTS U2033 ( .A(n2929), .B(n2930), .Y(n2918) );
  NOR2XLTS U2034 ( .A(n2942), .B(n2943), .Y(n2937) );
  NOR2XLTS U2035 ( .A(n2944), .B(n2743), .Y(n2943) );
  NOR2XLTS U2036 ( .A(n2763), .B(n2848), .Y(n2944) );
  NOR2XLTS U2037 ( .A(n2722), .B(n2947), .Y(n2942) );
  NOR2XLTS U2038 ( .A(n2948), .B(n2949), .Y(n2914) );
  NOR2XLTS U2039 ( .A(n3081), .B(n3082), .Y(n2951) );
  NOR2XLTS U2040 ( .A(n3086), .B(n3087), .Y(n3083) );
  NOR2XLTS U2041 ( .A(n3088), .B(n2829), .Y(n3086) );
  NOR2XLTS U2042 ( .A(n3093), .B(n3094), .Y(n3090) );
  NOR2XLTS U2043 ( .A(n3095), .B(n2813), .Y(n3094) );
  NOR2XLTS U2044 ( .A(n2778), .B(n2869), .Y(n3095) );
  NOR2XLTS U2045 ( .A(n3016), .B(n2740), .Y(n3093) );
  NOR2XLTS U2046 ( .A(n2816), .B(n2784), .Y(n3016) );
  NOR2XLTS U2047 ( .A(n2952), .B(n2953), .Y(n2950) );
  NOR2XLTS U2048 ( .A(n3146), .B(n3147), .Y(n3145) );
  NOR2XLTS U2049 ( .A(n3151), .B(n2803), .Y(n3146) );
  NOR2XLTS U2050 ( .A(n3152), .B(n3153), .Y(n3144) );
  NOR2XLTS U2051 ( .A(n2873), .B(n2859), .Y(n3158) );
  NOR2XLTS U2052 ( .A(n2750), .B(n2863), .Y(n2982) );
  NOR2XLTS U2053 ( .A(n2838), .B(n2802), .Y(n2952) );
  NOR2XLTS U2054 ( .A(n2957), .B(n2958), .Y(n2956) );
  NOR2XLTS U2055 ( .A(n3071), .B(n3072), .Y(n2959) );
  NOR2XLTS U2056 ( .A(n3078), .B(n3079), .Y(n3075) );
  NOR2XLTS U2057 ( .A(n2715), .B(n2776), .Y(n3079) );
  NOR2XLTS U2058 ( .A(n2757), .B(n2826), .Y(n3078) );
  NOR2XLTS U2059 ( .A(n3247), .B(n3508), .Y(n3164) );
  OR2XLTS U2060 ( .A(n3057), .B(n3509), .Y(n3508) );
  NOR2XLTS U2061 ( .A(n3512), .B(n3513), .Y(n3511) );
  NOR2XLTS U2062 ( .A(n3516), .B(n3517), .Y(n3514) );
  NOR2XLTS U2063 ( .A(n3187), .B(n2772), .Y(n3517) );
  NOR2XLTS U2064 ( .A(n3518), .B(n2768), .Y(n3516) );
  NOR2XLTS U2065 ( .A(n2842), .B(n2786), .Y(n3518) );
  NOR2XLTS U2066 ( .A(n3218), .B(n2752), .Y(n3512) );
  NOR2XLTS U2067 ( .A(n3519), .B(n3520), .Y(n3510) );
  INVXLTS U2068 ( .A(n3222), .Y(n3458) );
  NOR2XLTS U2069 ( .A(n3525), .B(n2828), .Y(n3519) );
  NOR2XLTS U2070 ( .A(n2702), .B(n3136), .Y(n3525) );
  NOR2XLTS U2071 ( .A(n3530), .B(n3531), .Y(n3529) );
  NOR2XLTS U2072 ( .A(n3151), .B(n2736), .Y(n3531) );
  NOR2XLTS U2073 ( .A(n3532), .B(n2732), .Y(n3530) );
  NOR2XLTS U2074 ( .A(n2875), .B(n3424), .Y(n3532) );
  NOR2XLTS U2075 ( .A(n3533), .B(n3534), .Y(n3528) );
  NOR2XLTS U2076 ( .A(n3536), .B(n3537), .Y(n3535) );
  NOR2XLTS U2077 ( .A(n2704), .B(n2802), .Y(n3537) );
  NOR2XLTS U2078 ( .A(n3169), .B(n2834), .Y(n3536) );
  NOR2XLTS U2079 ( .A(n3110), .B(n2807), .Y(n3533) );
  INVXLTS U2080 ( .A(n3136), .Y(n3110) );
  NOR2XLTS U2081 ( .A(n2740), .B(n2723), .Y(n3172) );
  NOR2XLTS U2082 ( .A(n3175), .B(n3176), .Y(n3174) );
  NOR2XLTS U2083 ( .A(n3432), .B(n3433), .Y(n3430) );
  NOR2XLTS U2084 ( .A(n3179), .B(n3180), .Y(n3178) );
  INVXLTS U2085 ( .A(n3184), .Y(n3183) );
  NOR2XLTS U2086 ( .A(n3185), .B(n3186), .Y(n3181) );
  NOR2XLTS U2087 ( .A(n3187), .B(n2826), .Y(n3186) );
  NOR2XLTS U2088 ( .A(n2873), .B(n2877), .Y(n3187) );
  NOR2XLTS U2089 ( .A(n3188), .B(n2813), .Y(n3185) );
  NOR2XLTS U2090 ( .A(n2887), .B(n2879), .Y(n3188) );
  NOR2XLTS U2091 ( .A(n3189), .B(n3190), .Y(n3177) );
  NOR2XLTS U2092 ( .A(n3195), .B(n2705), .Y(n3189) );
  NOR2XLTS U2093 ( .A(n2845), .B(n2934), .Y(n3195) );
  NOR2XLTS U2094 ( .A(n3196), .B(n3197), .Y(n3173) );
  NOR2XLTS U2095 ( .A(n3200), .B(n3201), .Y(n3198) );
  NOR2XLTS U2096 ( .A(n2819), .B(n2835), .Y(n3201) );
  NOR2XLTS U2097 ( .A(n2801), .B(n2752), .Y(n3200) );
  NOR2XLTS U2098 ( .A(n3087), .B(n3206), .Y(n3205) );
  NOR2XLTS U2099 ( .A(n2830), .B(n2742), .Y(n3206) );
  NOR2XLTS U2100 ( .A(n2760), .B(n2721), .Y(n3087) );
  NOR2XLTS U2101 ( .A(n3207), .B(n3208), .Y(n3204) );
  NOR2XLTS U2102 ( .A(n3015), .B(n2827), .Y(n3208) );
  NOR2XLTS U2103 ( .A(n3104), .B(n2789), .Y(n3207) );
  NOR2XLTS U2104 ( .A(n3211), .B(n3212), .Y(n3210) );
  NOR2XLTS U2105 ( .A(n3184), .B(n2835), .Y(n3212) );
  NOR2XLTS U2106 ( .A(n2764), .B(n2841), .Y(n3184) );
  NOR2XLTS U2107 ( .A(n3213), .B(n2795), .Y(n3211) );
  NOR2XLTS U2108 ( .A(n2933), .B(n3166), .Y(n3213) );
  NOR2XLTS U2109 ( .A(n3214), .B(n3215), .Y(n3209) );
  NOR2XLTS U2110 ( .A(n3218), .B(n2807), .Y(n3214) );
  NOR2XLTS U2111 ( .A(n2779), .B(n2882), .Y(n3218) );
  NOR2XLTS U2112 ( .A(n3364), .B(n3489), .Y(n3488) );
  NOR2XLTS U2113 ( .A(n3492), .B(n3493), .Y(n3490) );
  NOR2XLTS U2114 ( .A(n2829), .B(n2722), .Y(n3493) );
  NOR2XLTS U2115 ( .A(n2780), .B(n2792), .Y(n3492) );
  NOR2XLTS U2116 ( .A(n3494), .B(n3495), .Y(n3487) );
  NOR2XLTS U2117 ( .A(n2717), .B(n2756), .Y(n3498) );
  NOR2XLTS U2118 ( .A(n2769), .B(n2849), .Y(n3047) );
  NOR2XLTS U2119 ( .A(n3504), .B(n3505), .Y(n3501) );
  NOR2XLTS U2120 ( .A(n3506), .B(n2753), .Y(n3505) );
  NOR2XLTS U2121 ( .A(n2878), .B(n2744), .Y(n3506) );
  NOR2XLTS U2122 ( .A(n3507), .B(n2724), .Y(n3504) );
  NOR2XLTS U2123 ( .A(n2883), .B(n2725), .Y(n3507) );
  NOR2XLTS U2124 ( .A(n3225), .B(n2715), .Y(n3224) );
  NOR2XLTS U2125 ( .A(n2809), .B(n2934), .Y(n3225) );
  NOR2XLTS U2126 ( .A(n2813), .B(n3167), .Y(n3223) );
  NOR2XLTS U2127 ( .A(n3226), .B(n3227), .Y(n3031) );
  NOR2XLTS U2128 ( .A(n3230), .B(n3231), .Y(n3228) );
  NOR2XLTS U2129 ( .A(n2881), .B(n2860), .Y(n3088) );
  NOR2XLTS U2130 ( .A(n3235), .B(n2796), .Y(n3230) );
  NOR2XLTS U2131 ( .A(n2879), .B(n2747), .Y(n3235) );
  NOR2XLTS U2132 ( .A(n3238), .B(n3239), .Y(n3237) );
  AND2XLTS U2133 ( .A(n3244), .B(n3245), .Y(n3242) );
  INVXLTS U2134 ( .A(n2839), .Y(n3004) );
  NOR2XLTS U2135 ( .A(n3123), .B(n3246), .Y(n3236) );
  NOR2XLTS U2136 ( .A(n3109), .B(n2734), .Y(n3246) );
  NOR2XLTS U2137 ( .A(n3202), .B(n2828), .Y(n3123) );
  NOR2XLTS U2138 ( .A(n3438), .B(n3439), .Y(n3248) );
  OR2XLTS U2139 ( .A(n3440), .B(n3441), .Y(n3439) );
  NOR2XLTS U2140 ( .A(n3450), .B(n3451), .Y(n3449) );
  NOR2XLTS U2141 ( .A(n3222), .B(n2733), .Y(n3451) );
  NOR2XLTS U2142 ( .A(n3171), .B(n2793), .Y(n3450) );
  NOR2XLTS U2143 ( .A(n3452), .B(n3453), .Y(n3448) );
  NOR2XLTS U2144 ( .A(n3456), .B(n3457), .Y(n3454) );
  NOR2XLTS U2145 ( .A(n2796), .B(n2835), .Y(n3457) );
  NOR2XLTS U2146 ( .A(n2767), .B(n2814), .Y(n3456) );
  NOR2XLTS U2147 ( .A(n2941), .B(n2824), .Y(n3452) );
  NOR2XLTS U2148 ( .A(n2852), .B(n2855), .Y(n2941) );
  NOR2XLTS U2149 ( .A(n3251), .B(n3252), .Y(n3250) );
  NOR2XLTS U2150 ( .A(n3259), .B(n3260), .Y(n3249) );
  NOR2XLTS U2151 ( .A(n3059), .B(n3540), .Y(n3539) );
  NOR2XLTS U2152 ( .A(n3545), .B(n3546), .Y(n3541) );
  INVXLTS U2153 ( .A(n3134), .Y(n3040) );
  NOR2XLTS U2154 ( .A(n2873), .B(n2779), .Y(n3544) );
  NOR2XLTS U2155 ( .A(n3564), .B(n3565), .Y(n3557) );
  NOR2XLTS U2156 ( .A(n3572), .B(n2757), .Y(n3564) );
  NOR2XLTS U2157 ( .A(n2810), .B(n3574), .Y(n3572) );
  NOR2XLTS U2158 ( .A(n3058), .B(n3575), .Y(n3538) );
  NOR2XLTS U2159 ( .A(n3411), .B(n3582), .Y(n3581) );
  NOR2XLTS U2160 ( .A(n2822), .B(n2771), .Y(n3582) );
  NOR2XLTS U2161 ( .A(n3584), .B(n3585), .Y(n3580) );
  NOR2XLTS U2162 ( .A(n3171), .B(n2805), .Y(n3585) );
  NOR2XLTS U2163 ( .A(n2858), .B(n2745), .Y(n3171) );
  NOR2XLTS U2164 ( .A(n3588), .B(n2720), .Y(n3584) );
  NOR2XLTS U2165 ( .A(n2817), .B(n2854), .Y(n3588) );
  NOR2XLTS U2166 ( .A(n3270), .B(n3271), .Y(n3269) );
  NOR2XLTS U2167 ( .A(n2957), .B(n2968), .Y(n3273) );
  NOR2XLTS U2168 ( .A(n3276), .B(n3277), .Y(n3275) );
  NOR2XLTS U2169 ( .A(n3282), .B(n3036), .Y(n3280) );
  NOR2XLTS U2170 ( .A(n2800), .B(n2814), .Y(n3036) );
  NOR2XLTS U2171 ( .A(n2826), .B(n2742), .Y(n3282) );
  NOR2XLTS U2172 ( .A(n3283), .B(n3284), .Y(n3274) );
  INVXLTS U2173 ( .A(n3288), .Y(n3104) );
  NOR2XLTS U2174 ( .A(n2912), .B(n3289), .Y(n3132) );
  NOR2XLTS U2175 ( .A(n3293), .B(n3294), .Y(n3290) );
  NOR2XLTS U2176 ( .A(n3109), .B(n2766), .Y(n3294) );
  NOR2XLTS U2177 ( .A(n2717), .B(n2738), .Y(n3109) );
  NOR2XLTS U2178 ( .A(n3295), .B(n2861), .Y(n3293) );
  NOR2XLTS U2179 ( .A(n3298), .B(n3299), .Y(n3297) );
  NOR2XLTS U2180 ( .A(n2954), .B(n2831), .Y(n3299) );
  NOR2XLTS U2181 ( .A(n2806), .B(n2822), .Y(n3298) );
  NOR2XLTS U2182 ( .A(n3300), .B(n3301), .Y(n3296) );
  NOR2XLTS U2183 ( .A(n2794), .B(n2710), .Y(n3300) );
  NOR2XLTS U2184 ( .A(n3305), .B(n3306), .Y(n3272) );
  NOR2XLTS U2185 ( .A(n3309), .B(n3310), .Y(n3308) );
  NOR2XLTS U2186 ( .A(n2716), .B(n2805), .Y(n3310) );
  NOR2XLTS U2187 ( .A(n2710), .B(n2827), .Y(n3309) );
  NOR2XLTS U2188 ( .A(n3311), .B(n3312), .Y(n3307) );
  NOR2XLTS U2189 ( .A(n2720), .B(n2815), .Y(n3312) );
  NOR2XLTS U2190 ( .A(n3151), .B(n2775), .Y(n3311) );
  NOR2XLTS U2191 ( .A(n2730), .B(n3085), .Y(n3151) );
  NOR2XLTS U2192 ( .A(n3315), .B(n3316), .Y(n3314) );
  NOR2XLTS U2193 ( .A(n3014), .B(n2833), .Y(n3316) );
  NOR2XLTS U2194 ( .A(n2693), .B(n2765), .Y(n3014) );
  NOR2XLTS U2195 ( .A(n3317), .B(n2790), .Y(n3315) );
  NOR2XLTS U2196 ( .A(n2701), .B(n3257), .Y(n3317) );
  NOR2XLTS U2197 ( .A(n3318), .B(n3319), .Y(n3313) );
  NOR2XLTS U2198 ( .A(n3320), .B(n2727), .Y(n3319) );
  NOR2XLTS U2199 ( .A(n2844), .B(n2851), .Y(n3320) );
  NOR2XLTS U2200 ( .A(n3321), .B(n2800), .Y(n3318) );
  NOR2XLTS U2201 ( .A(n2783), .B(n2809), .Y(n3321) );
  OR2XLTS U2202 ( .A(n3019), .B(n3322), .Y(n3270) );
  NOR2XLTS U2203 ( .A(n3324), .B(n3325), .Y(n3323) );
  NOR2XLTS U2204 ( .A(n2762), .B(n2742), .Y(n3325) );
  NOR2XLTS U2205 ( .A(n2820), .B(n2759), .Y(n3324) );
  NOR2XLTS U2206 ( .A(n3326), .B(n3327), .Y(n2960) );
  NOR2XLTS U2207 ( .A(n2798), .B(n2738), .Y(n2977) );
  NOR2XLTS U2208 ( .A(n3334), .B(n3335), .Y(n3331) );
  NOR2XLTS U2209 ( .A(n3336), .B(n2793), .Y(n3335) );
  NOR2XLTS U2210 ( .A(n2882), .B(n2870), .Y(n3336) );
  NOR2XLTS U2211 ( .A(n3337), .B(n2834), .Y(n3334) );
  NOR2XLTS U2212 ( .A(n2718), .B(n2816), .Y(n3337) );
  NOR2XLTS U2213 ( .A(n3340), .B(n3341), .Y(n3339) );
  INVXLTS U2214 ( .A(n2740), .Y(n3023) );
  NOR2XLTS U2215 ( .A(n3345), .B(n3346), .Y(n3338) );
  NOR2XLTS U2216 ( .A(n2871), .B(n2859), .Y(n3350) );
  NOR2XLTS U2217 ( .A(n2695), .B(n2713), .Y(n3169) );
  INVXLTS U2218 ( .A(n2792), .Y(n3097) );
  INVXLTS U2219 ( .A(n2795), .Y(n2924) );
  NOR2XLTS U2220 ( .A(n2797), .B(n2842), .Y(n3295) );
  NOR2XLTS U2221 ( .A(n3523), .B(n3289), .Y(n2986) );
  NOR2XLTS U2222 ( .A(n2811), .B(n2714), .Y(n3222) );
  NOR2XLTS U2223 ( .A(n3568), .B(n3573), .Y(n2928) );
  NOR2XLTS U2224 ( .A(n3363), .B(n2788), .Y(n3357) );
  NOR2XLTS U2225 ( .A(n2869), .B(n2696), .Y(n3363) );
  INVXLTS U2226 ( .A(n2824), .Y(n3006) );
  NOR2XLTS U2227 ( .A(n3364), .B(n3365), .Y(n3017) );
  NOR2XLTS U2228 ( .A(n3368), .B(n3369), .Y(n3366) );
  NOR2XLTS U2229 ( .A(n2830), .B(n2710), .Y(n3369) );
  NOR2XLTS U2230 ( .A(n2803), .B(n3167), .Y(n3368) );
  NOR2XLTS U2231 ( .A(n2821), .B(n2823), .Y(n3364) );
  NOR2XLTS U2232 ( .A(n3371), .B(n3372), .Y(n2955) );
  NOR2XLTS U2233 ( .A(n3375), .B(n3376), .Y(n3374) );
  NOR2XLTS U2234 ( .A(n2835), .B(n2731), .Y(n3376) );
  NOR2XLTS U2235 ( .A(n2739), .B(n2752), .Y(n3375) );
  NOR2XLTS U2236 ( .A(n3377), .B(n3378), .Y(n3373) );
  NOR2XLTS U2237 ( .A(n2733), .B(n2789), .Y(n3377) );
  NOR2XLTS U2238 ( .A(n3382), .B(n3383), .Y(n3381) );
  NOR2XLTS U2239 ( .A(n2711), .B(n2762), .Y(n3383) );
  NOR2XLTS U2240 ( .A(n3384), .B(n2791), .Y(n3382) );
  NOR2XLTS U2241 ( .A(n2886), .B(n2862), .Y(n3384) );
  NOR2XLTS U2242 ( .A(n3385), .B(n3386), .Y(n3380) );
  NOR2XLTS U2243 ( .A(n3390), .B(n2820), .Y(n3385) );
  NOR2XLTS U2244 ( .A(n2729), .B(n3115), .Y(n3390) );
  NOR2XLTS U2245 ( .A(n3392), .B(n3393), .Y(n3018) );
  NOR2XLTS U2246 ( .A(n2909), .B(n2912), .Y(n3561) );
  INVXLTS U2247 ( .A(n2734), .Y(n3085) );
  NOR2XLTS U2248 ( .A(n3402), .B(n3403), .Y(n3399) );
  NOR2XLTS U2249 ( .A(n3404), .B(n2761), .Y(n3403) );
  NOR2XLTS U2250 ( .A(n3405), .B(n2728), .Y(n3402) );
  NOR2XLTS U2251 ( .A(n2841), .B(n2737), .Y(n3405) );
  NOR2XLTS U2252 ( .A(n3406), .B(n3407), .Y(n2965) );
  NOR2XLTS U2253 ( .A(n3410), .B(n3411), .Y(n3409) );
  NOR2XLTS U2254 ( .A(n2802), .B(n2834), .Y(n3411) );
  NOR2XLTS U2255 ( .A(n2723), .B(n2733), .Y(n3410) );
  NOR2XLTS U2256 ( .A(n3412), .B(n3413), .Y(n3408) );
  NOR2XLTS U2257 ( .A(n2731), .B(n2823), .Y(n3413) );
  INVXLTS U2258 ( .A(n3398), .Y(n3304) );
  NOR2XLTS U2259 ( .A(n2727), .B(n2814), .Y(n3412) );
  NOR2XLTS U2260 ( .A(n3416), .B(n3417), .Y(n3415) );
  NOR2XLTS U2261 ( .A(n3418), .B(n2772), .Y(n3417) );
  NOR2XLTS U2262 ( .A(n3461), .B(n3583), .Y(n3051) );
  INVXLTS U2263 ( .A(n3499), .Y(n3461) );
  NOR2XLTS U2264 ( .A(n2857), .B(n3288), .Y(n3418) );
  NOR2XLTS U2265 ( .A(n3523), .B(n3524), .Y(n2975) );
  NOR2XLTS U2266 ( .A(n3556), .B(n3289), .Y(n2939) );
  NOR2XLTS U2267 ( .A(n3419), .B(n2806), .Y(n3416) );
  NOR2XLTS U2268 ( .A(n2903), .B(n3398), .Y(n2946) );
  NOR2XLTS U2269 ( .A(n2874), .B(n2862), .Y(n3419) );
  NOR2XLTS U2270 ( .A(n3526), .B(n3527), .Y(n2933) );
  NOR2XLTS U2271 ( .A(n3523), .B(n3563), .Y(n2994) );
  OR2XLTS U2272 ( .A(n2891), .B(n2908), .Y(n3563) );
  INVXLTS U2273 ( .A(n3466), .Y(n3523) );
  NOR2XLTS U2274 ( .A(n3420), .B(n3421), .Y(n3414) );
  NOR2XLTS U2275 ( .A(n3556), .B(n3524), .Y(n2925) );
  NOR2XLTS U2276 ( .A(n3526), .B(n3556), .Y(n3077) );
  INVXLTS U2277 ( .A(n2729), .Y(n3015) );
  NOR2XLTS U2278 ( .A(n2708), .B(n3583), .Y(n3161) );
  INVXLTS U2279 ( .A(n3586), .Y(n3583) );
  NOR2XLTS U2280 ( .A(n2893), .B(n2906), .Y(n3586) );
  NOR2XLTS U2281 ( .A(n3426), .B(n3427), .Y(n3420) );
  AND2XLTS U2282 ( .A(n2899), .B(n2902), .Y(n3428) );
  NOR2XLTS U2283 ( .A(n2911), .B(n3570), .Y(n3587) );
  INVXLTS U2284 ( .A(n3568), .Y(n3560) );
  OR2XLTS U2285 ( .A(n2896), .B(n2891), .Y(n3568) );
  NOR2XLTS U2286 ( .A(n2896), .B(n3289), .Y(n3446) );
  INVXLTS U2287 ( .A(n2908), .Y(n3570) );
  NOR2XLTS U2288 ( .A(n3526), .B(n3578), .Y(n2935) );
  INVXLTS U2289 ( .A(n2911), .Y(n3562) );
  INVXLTS U2290 ( .A(n3370), .Y(n3526) );
  AND2XLTS U2291 ( .A(n2890), .B(n2909), .Y(n3370) );
  NOR2XLTS U2292 ( .A(n3004), .B(n2875), .Y(n3003) );
  NOR2XLTS U2293 ( .A(n2866), .B(n2883), .Y(n3404) );
  NAND2X1TS U2294 ( .A(n3499), .B(n3500), .Y(n3131) );
  NOR2BX1TS U2295 ( .AN(n2906), .B(n2894), .Y(n3500) );
  NOR2X1TS U2296 ( .A(n2902), .B(n2900), .Y(n3499) );
  NOR2BX1TS U2297 ( .AN(n2897), .B(n2913), .Y(n3466) );
  NOR2BX1TS U2298 ( .AN(n2894), .B(n2905), .Y(n3459) );
  NOR2BX1TS U2299 ( .AN(n2900), .B(n2902), .Y(n3555) );
  NAND2X1TS U2300 ( .A(n2912), .B(n2896), .Y(n3556) );
  NOR2BX1TS U2301 ( .AN(n2903), .B(n2899), .Y(n3460) );
  NAND2X1TS U2302 ( .A(n2890), .B(n3570), .Y(n3289) );
  NAND2X1TS U2303 ( .A(n3466), .B(n2889), .Y(n3465) );
  NAND2X1TS U2304 ( .A(n2961), .B(n2962), .Y(d[6]) );
  NAND2X1TS U2305 ( .A(n2965), .B(n2966), .Y(n2964) );
  NAND2X1TS U2306 ( .A(n2969), .B(n2970), .Y(n2967) );
  NAND2X1TS U2307 ( .A(n2973), .B(n2974), .Y(n2972) );
  NAND2X1TS U2308 ( .A(n2870), .B(n2738), .Y(n2974) );
  NAND2X1TS U2309 ( .A(n2817), .B(n2976), .Y(n2973) );
  NAND2X1TS U2310 ( .A(n2980), .B(n2981), .Y(n2979) );
  NAND2BX1TS U2311 ( .AN(n2982), .B(n2810), .Y(n2981) );
  NAND2X1TS U2312 ( .A(n2786), .B(n2983), .Y(n2980) );
  NAND2X1TS U2313 ( .A(n2780), .B(n2758), .Y(n2983) );
  NAND2X1TS U2314 ( .A(n2984), .B(n2985), .Y(n2978) );
  NAND2X1TS U2315 ( .A(n2859), .B(n2987), .Y(n2985) );
  NAND2X1TS U2316 ( .A(n2791), .B(n2753), .Y(n2987) );
  NAND2X1TS U2317 ( .A(n2844), .B(n2989), .Y(n2984) );
  NAND2X1TS U2318 ( .A(n2990), .B(n2823), .Y(n2989) );
  NAND2X1TS U2319 ( .A(n2992), .B(n2993), .Y(n2991) );
  NAND2X1TS U2320 ( .A(n2718), .B(n2883), .Y(n2993) );
  NAND2X1TS U2321 ( .A(n2994), .B(n2769), .Y(n2992) );
  NAND2X1TS U2322 ( .A(n3026), .B(n3027), .Y(d[5]) );
  NAND2X1TS U2323 ( .A(n3030), .B(n3031), .Y(n3029) );
  NAND2X1TS U2324 ( .A(n3034), .B(n3035), .Y(n3033) );
  NAND2X1TS U2325 ( .A(n3041), .B(n3042), .Y(n3032) );
  NAND2X1TS U2326 ( .A(n2727), .B(n3045), .Y(n2976) );
  NAND2X1TS U2327 ( .A(n2908), .B(n3046), .Y(n3045) );
  NAND2X1TS U2328 ( .A(n3468), .B(n3469), .Y(n3467) );
  NAND2X1TS U2329 ( .A(n3472), .B(n3473), .Y(n3471) );
  NAND2X1TS U2330 ( .A(n2873), .B(n2751), .Y(n3473) );
  NAND2X1TS U2331 ( .A(n2852), .B(n3424), .Y(n3472) );
  NAND2X1TS U2332 ( .A(n3476), .B(n3477), .Y(n3475) );
  NAND2X1TS U2333 ( .A(n3051), .B(n3156), .Y(n3477) );
  NAND2X1TS U2334 ( .A(n2810), .B(n3478), .Y(n3476) );
  NAND2X1TS U2335 ( .A(n2834), .B(n2768), .Y(n3478) );
  NAND2X1TS U2336 ( .A(n3479), .B(n3480), .Y(n3474) );
  NAND2X1TS U2337 ( .A(n2870), .B(n3481), .Y(n3480) );
  NAND2X1TS U2338 ( .A(n2827), .B(n3482), .Y(n3481) );
  NAND2X1TS U2339 ( .A(n2906), .B(n2709), .Y(n3482) );
  NAND2X1TS U2340 ( .A(n3054), .B(n3055), .Y(n3052) );
  NAND2X1TS U2341 ( .A(n3060), .B(n3061), .Y(d[4]) );
  NAND2X1TS U2342 ( .A(n3063), .B(n3064), .Y(n3062) );
  NOR2BX1TS U2343 ( .AN(n2951), .B(n3065), .Y(n3064) );
  NAND2X1TS U2344 ( .A(n2959), .B(n3066), .Y(n3065) );
  NAND2X1TS U2345 ( .A(n3069), .B(n3070), .Y(n3068) );
  NAND2X1TS U2346 ( .A(n2845), .B(n2859), .Y(n3069) );
  NAND2X1TS U2347 ( .A(n3100), .B(n3101), .Y(n3099) );
  NAND2X1TS U2348 ( .A(n2747), .B(n3102), .Y(n3101) );
  NAND2X1TS U2349 ( .A(n2760), .B(n2826), .Y(n3102) );
  NAND2X1TS U2350 ( .A(n2754), .B(n3103), .Y(n3100) );
  NAND2X1TS U2351 ( .A(n3104), .B(n2758), .Y(n3103) );
  NAND2X1TS U2352 ( .A(n3105), .B(n3106), .Y(n3098) );
  NAND2X1TS U2353 ( .A(n3113), .B(n3114), .Y(n3112) );
  NAND2X1TS U2354 ( .A(n2726), .B(n2786), .Y(n3114) );
  NAND2X1TS U2355 ( .A(n2769), .B(n3115), .Y(n3113) );
  NAND2X1TS U2356 ( .A(n3117), .B(n3118), .Y(n3116) );
  NAND2X1TS U2357 ( .A(n3121), .B(n3122), .Y(n3120) );
  NAND2X1TS U2358 ( .A(n3128), .B(n3129), .Y(n3127) );
  NAND2X1TS U2359 ( .A(n2871), .B(n3130), .Y(n3129) );
  NAND2X1TS U2360 ( .A(n2821), .B(n2724), .Y(n3130) );
  NAND2X1TS U2361 ( .A(n2770), .B(n3132), .Y(n3128) );
  NAND2X1TS U2362 ( .A(n3139), .B(n3140), .Y(n3138) );
  NAND2X1TS U2363 ( .A(n2862), .B(n2852), .Y(n3140) );
  NAND2X1TS U2364 ( .A(n2748), .B(n2785), .Y(n3139) );
  NAND2X1TS U2365 ( .A(n3142), .B(n3143), .Y(n3137) );
  NAND2X1TS U2366 ( .A(n2755), .B(n2779), .Y(n3143) );
  NAND2X1TS U2367 ( .A(n2865), .B(n2848), .Y(n3142) );
  NAND2X1TS U2368 ( .A(n2914), .B(n2915), .Y(d[7]) );
  NAND2X1TS U2369 ( .A(n2995), .B(n2996), .Y(n2917) );
  NAND2X1TS U2370 ( .A(n2999), .B(n3000), .Y(n2998) );
  NAND2X1TS U2371 ( .A(n3009), .B(n3010), .Y(n3008) );
  NAND2X1TS U2372 ( .A(n2725), .B(n2713), .Y(n3010) );
  NAND2X1TS U2373 ( .A(n3017), .B(n3018), .Y(n2997) );
  NAND2X1TS U2374 ( .A(n3021), .B(n3022), .Y(n3020) );
  NAND2X1TS U2375 ( .A(n2750), .B(n2755), .Y(n3022) );
  NAND2X1TS U2376 ( .A(n2918), .B(n2919), .Y(n2916) );
  NAND2X1TS U2377 ( .A(n2922), .B(n2923), .Y(n2921) );
  NAND2X1TS U2378 ( .A(n2729), .B(n2817), .Y(n2923) );
  NAND2X1TS U2379 ( .A(n2882), .B(n2797), .Y(n2922) );
  NAND2X1TS U2380 ( .A(n2926), .B(n2927), .Y(n2920) );
  NAND2X1TS U2381 ( .A(n2770), .B(n2878), .Y(n2927) );
  NAND2X1TS U2382 ( .A(n2811), .B(n2702), .Y(n2926) );
  NAND2X1TS U2383 ( .A(n2931), .B(n2932), .Y(n2930) );
  NAND2X1TS U2384 ( .A(n2863), .B(n2934), .Y(n2932) );
  NAND2X1TS U2385 ( .A(n2887), .B(n2936), .Y(n2931) );
  NAND2X1TS U2386 ( .A(n2937), .B(n2938), .Y(n2929) );
  NAND2X1TS U2387 ( .A(n2857), .B(n2940), .Y(n2938) );
  NAND2X1TS U2388 ( .A(n2941), .B(n2791), .Y(n2940) );
  NAND2X1TS U2389 ( .A(n2706), .B(n2898), .Y(n2947) );
  NAND2X1TS U2390 ( .A(n2950), .B(n2951), .Y(n2949) );
  NAND2X1TS U2391 ( .A(n3083), .B(n3084), .Y(n3082) );
  NAND2X1TS U2392 ( .A(n2816), .B(n2778), .Y(n3084) );
  NAND2X1TS U2393 ( .A(n3090), .B(n3091), .Y(n3081) );
  NAND2X1TS U2394 ( .A(n2845), .B(n3092), .Y(n3091) );
  NAND2X1TS U2395 ( .A(n2712), .B(n2720), .Y(n3092) );
  NAND2X1TS U2396 ( .A(n3144), .B(n3145), .Y(n2953) );
  NAND2X1TS U2397 ( .A(n3148), .B(n3149), .Y(n3147) );
  NAND2X1TS U2398 ( .A(n2875), .B(n3150), .Y(n3149) );
  NAND2X1TS U2399 ( .A(n2811), .B(n2745), .Y(n3148) );
  NAND2X1TS U2400 ( .A(n3154), .B(n3155), .Y(n3153) );
  NAND2X1TS U2401 ( .A(n2784), .B(n3156), .Y(n3155) );
  NAND2X1TS U2402 ( .A(n2954), .B(n2781), .Y(n3156) );
  NAND2X1TS U2403 ( .A(n2787), .B(n3157), .Y(n3154) );
  NAND2X1TS U2404 ( .A(n3158), .B(n2727), .Y(n3157) );
  NAND2X1TS U2405 ( .A(n3159), .B(n3160), .Y(n3152) );
  NAND2X1TS U2406 ( .A(n2855), .B(n3162), .Y(n3160) );
  NAND2X1TS U2407 ( .A(n2982), .B(n2721), .Y(n3162) );
  NAND2X1TS U2408 ( .A(n2879), .B(n3163), .Y(n3159) );
  NAND2X1TS U2409 ( .A(n2796), .B(n2789), .Y(n3163) );
  NAND2X1TS U2410 ( .A(n2955), .B(n2956), .Y(n2948) );
  NAND2X1TS U2411 ( .A(n2959), .B(n2960), .Y(n2958) );
  NAND2X1TS U2412 ( .A(n3073), .B(n3074), .Y(n3072) );
  NAND2X1TS U2413 ( .A(n2885), .B(n2849), .Y(n3074) );
  NAND2X1TS U2414 ( .A(n2798), .B(n2725), .Y(n3073) );
  NAND2X1TS U2415 ( .A(n3075), .B(n3076), .Y(n3071) );
  NAND2X1TS U2416 ( .A(n2865), .B(n2842), .Y(n3076) );
  NAND2X1TS U2417 ( .A(n3510), .B(n3511), .Y(n3509) );
  NAND2X1TS U2418 ( .A(n3514), .B(n3515), .Y(n3513) );
  NAND2X1TS U2419 ( .A(n2855), .B(n3257), .Y(n3515) );
  NAND2X1TS U2420 ( .A(n3521), .B(n3522), .Y(n3520) );
  NAND2X1TS U2421 ( .A(n2816), .B(n2874), .Y(n3522) );
  NAND2X1TS U2422 ( .A(n2869), .B(n3458), .Y(n3521) );
  NAND2X1TS U2423 ( .A(n3528), .B(n3529), .Y(n3057) );
  NAND2X1TS U2424 ( .A(n3535), .B(n3342), .Y(n3534) );
  NAND2X1TS U2425 ( .A(n2766), .B(n2822), .Y(n3136) );
  NAND2X1TS U2426 ( .A(n3169), .B(n2788), .Y(n3168) );
  NAND2X1TS U2427 ( .A(n2753), .B(n2736), .Y(n3170) );
  NAND2X1TS U2428 ( .A(n2717), .B(n2887), .Y(n3070) );
  NAND2X1TS U2429 ( .A(n3173), .B(n3174), .Y(n3028) );
  NAND2X1TS U2430 ( .A(n3430), .B(n3431), .Y(n3176) );
  NAND2X1TS U2431 ( .A(n2747), .B(n2713), .Y(n3431) );
  NAND2X1TS U2432 ( .A(n3434), .B(n3435), .Y(n3433) );
  NAND2X1TS U2433 ( .A(n2863), .B(n2787), .Y(n3435) );
  NAND2X1TS U2434 ( .A(n2797), .B(n2860), .Y(n3434) );
  NAND2X1TS U2435 ( .A(n3436), .B(n3437), .Y(n3432) );
  NAND2X1TS U2436 ( .A(n2924), .B(n2866), .Y(n3437) );
  NAND2X1TS U2437 ( .A(n2754), .B(n2882), .Y(n3436) );
  NAND2X1TS U2438 ( .A(n3177), .B(n3178), .Y(n3175) );
  NAND2X1TS U2439 ( .A(n3181), .B(n3182), .Y(n3180) );
  NAND2X1TS U2440 ( .A(n2885), .B(n3183), .Y(n3182) );
  NAND2X1TS U2441 ( .A(n3191), .B(n3192), .Y(n3190) );
  NAND2X1TS U2442 ( .A(n2939), .B(n3193), .Y(n3192) );
  NAND2X1TS U2443 ( .A(n2795), .B(n2803), .Y(n3193) );
  NAND2X1TS U2444 ( .A(n2867), .B(n3194), .Y(n3191) );
  NAND2X1TS U2445 ( .A(n2820), .B(n2775), .Y(n3194) );
  NAND2X1TS U2446 ( .A(n3198), .B(n3199), .Y(n3197) );
  NAND2X1TS U2447 ( .A(n2849), .B(n2870), .Y(n3199) );
  NAND2X1TS U2448 ( .A(n3204), .B(n3205), .Y(n3179) );
  NAND2X1TS U2449 ( .A(n3209), .B(n3210), .Y(n3196) );
  NAND2X1TS U2450 ( .A(n2800), .B(n2743), .Y(n3166) );
  NAND2X1TS U2451 ( .A(n3216), .B(n3217), .Y(n3215) );
  NAND2BX1TS U2452 ( .AN(n2941), .B(n2860), .Y(n3217) );
  NAND2X1TS U2453 ( .A(n2854), .B(n3115), .Y(n3216) );
  NAND2X1TS U2454 ( .A(n3487), .B(n3488), .Y(n3203) );
  NAND2X1TS U2455 ( .A(n3490), .B(n3491), .Y(n3489) );
  NAND2X1TS U2456 ( .A(n2817), .B(n2886), .Y(n3491) );
  NAND2X1TS U2457 ( .A(n3496), .B(n3497), .Y(n3495) );
  NAND2X1TS U2458 ( .A(n3004), .B(n3150), .Y(n3497) );
  NAND2X1TS U2459 ( .A(n3498), .B(n2804), .Y(n3150) );
  NAND2BX1TS U2460 ( .AN(n3384), .B(n2852), .Y(n3496) );
  NAND2X1TS U2461 ( .A(n3501), .B(n3502), .Y(n3494) );
  NAND2X1TS U2462 ( .A(n2730), .B(n3503), .Y(n3502) );
  NAND2X1TS U2463 ( .A(n3047), .B(n2771), .Y(n3503) );
  NAND2X1TS U2464 ( .A(n2885), .B(n2783), .Y(n3220) );
  NAND2X1TS U2465 ( .A(n2755), .B(n2879), .Y(n3219) );
  NAND2X1TS U2466 ( .A(n3109), .B(n3222), .Y(n3221) );
  NAND2X1TS U2467 ( .A(n2790), .B(n2774), .Y(n2934) );
  NAND2X1TS U2468 ( .A(n3228), .B(n3229), .Y(n3227) );
  NAND2X1TS U2469 ( .A(n3006), .B(n2936), .Y(n3229) );
  NAND2X1TS U2470 ( .A(n2988), .B(n2731), .Y(n2936) );
  NAND2X1TS U2471 ( .A(n3232), .B(n3233), .Y(n3231) );
  NAND2BX1TS U2472 ( .AN(n3088), .B(n2765), .Y(n3233) );
  NAND2X1TS U2473 ( .A(n2844), .B(n3234), .Y(n3232) );
  NAND2X1TS U2474 ( .A(n2782), .B(n2716), .Y(n3234) );
  NAND2X1TS U2475 ( .A(n3236), .B(n3237), .Y(n3226) );
  NAND2X1TS U2476 ( .A(n3240), .B(n3241), .Y(n3239) );
  NAND2X1TS U2477 ( .A(n2729), .B(n2784), .Y(n3241) );
  NAND2X1TS U2478 ( .A(n3242), .B(n3243), .Y(n3238) );
  NAND2X1TS U2479 ( .A(n2888), .B(n2810), .Y(n3243) );
  NAND2X1TS U2480 ( .A(n3004), .B(n2770), .Y(n3245) );
  NAND2X1TS U2481 ( .A(n3442), .B(n3443), .Y(n3441) );
  NAND2X1TS U2482 ( .A(n2883), .B(n2737), .Y(n3443) );
  NAND2X1TS U2483 ( .A(n2770), .B(n3330), .Y(n3442) );
  NAND2X1TS U2484 ( .A(n3444), .B(n3445), .Y(n3440) );
  NAND2X1TS U2485 ( .A(n3446), .B(n2764), .Y(n3445) );
  NAND2X1TS U2486 ( .A(n2862), .B(n3447), .Y(n3444) );
  NAND2X1TS U2487 ( .A(n2819), .B(n2840), .Y(n3447) );
  NAND2X1TS U2488 ( .A(n3448), .B(n3449), .Y(n3438) );
  NAND2X1TS U2489 ( .A(n3454), .B(n3455), .Y(n3453) );
  NAND2X1TS U2490 ( .A(n2887), .B(n2785), .Y(n3455) );
  NAND2X1TS U2491 ( .A(n3249), .B(n3250), .Y(n3165) );
  NAND2X1TS U2492 ( .A(n3253), .B(n3254), .Y(n3252) );
  NAND2X1TS U2493 ( .A(n2750), .B(n2809), .Y(n3254) );
  NAND2X1TS U2494 ( .A(n2875), .B(n2714), .Y(n3253) );
  NAND2X1TS U2495 ( .A(n3255), .B(n3256), .Y(n3251) );
  NAND2X1TS U2496 ( .A(n2754), .B(n3257), .Y(n3256) );
  NAND2X1TS U2497 ( .A(n2860), .B(n3258), .Y(n3255) );
  NAND2X1TS U2498 ( .A(n3261), .B(n3262), .Y(n3260) );
  NAND2X1TS U2499 ( .A(n2763), .B(n3263), .Y(n3262) );
  NAND2X1TS U2500 ( .A(n3040), .B(n2782), .Y(n3263) );
  NAND2X1TS U2501 ( .A(n3006), .B(n3264), .Y(n3261) );
  NAND2X1TS U2502 ( .A(n2792), .B(n2776), .Y(n3264) );
  NAND2X1TS U2503 ( .A(n3265), .B(n3266), .Y(n3259) );
  NAND2X1TS U2504 ( .A(n2751), .B(n3267), .Y(n3266) );
  NAND2X1TS U2505 ( .A(n2711), .B(n2721), .Y(n3267) );
  NAND2X1TS U2506 ( .A(n2886), .B(n3268), .Y(n3265) );
  NAND2X1TS U2507 ( .A(n2805), .B(n2828), .Y(n3268) );
  NAND2X1TS U2508 ( .A(n3538), .B(n3539), .Y(n3247) );
  NAND2X1TS U2509 ( .A(n3541), .B(n3542), .Y(n3540) );
  NAND2X1TS U2510 ( .A(n2756), .B(n3543), .Y(n3542) );
  NAND2X1TS U2511 ( .A(n3544), .B(n2833), .Y(n3543) );
  NAND2X1TS U2512 ( .A(n3547), .B(n3548), .Y(n3546) );
  NAND2X1TS U2513 ( .A(n2783), .B(n3549), .Y(n3548) );
  NAND2X1TS U2514 ( .A(n2739), .B(n2767), .Y(n3549) );
  NAND2X1TS U2515 ( .A(n2846), .B(n3550), .Y(n3547) );
  NAND2X1TS U2516 ( .A(n3040), .B(n2733), .Y(n3550) );
  NAND2X1TS U2517 ( .A(n2839), .B(n2759), .Y(n3134) );
  NAND2X1TS U2518 ( .A(n3551), .B(n3552), .Y(n3545) );
  NAND2X1TS U2519 ( .A(n2925), .B(n3553), .Y(n3552) );
  NAND2X1TS U2520 ( .A(n3169), .B(n2775), .Y(n3553) );
  NAND2X1TS U2521 ( .A(n2866), .B(n3554), .Y(n3551) );
  NAND2X1TS U2522 ( .A(n2732), .B(n2827), .Y(n3554) );
  NAND2X1TS U2523 ( .A(n3557), .B(n3558), .Y(n3059) );
  NAND2X1TS U2524 ( .A(n3097), .B(n3559), .Y(n3558) );
  NAND2X1TS U2525 ( .A(n3544), .B(n2839), .Y(n3559) );
  NAND2X1TS U2526 ( .A(n3566), .B(n3567), .Y(n3565) );
  NAND2X1TS U2527 ( .A(n2756), .B(n3464), .Y(n3567) );
  NAND2X1TS U2528 ( .A(n3015), .B(n2766), .Y(n3464) );
  NAND2X1TS U2529 ( .A(n3023), .B(n3571), .Y(n3566) );
  NAND2X1TS U2530 ( .A(n2803), .B(n2752), .Y(n3571) );
  NAND2X1TS U2531 ( .A(n2774), .B(n2735), .Y(n3574) );
  NAND2X1TS U2532 ( .A(n3576), .B(n3577), .Y(n3575) );
  NAND2X1TS U2533 ( .A(n2888), .B(n2797), .Y(n3577) );
  NAND2X1TS U2534 ( .A(n2858), .B(n3579), .Y(n3576) );
  NAND2X1TS U2535 ( .A(n2761), .B(n2814), .Y(n3579) );
  NAND2X1TS U2536 ( .A(n3580), .B(n3581), .Y(n3058) );
  NAND2X1TS U2537 ( .A(n3060), .B(n3269), .Y(d[1]) );
  NAND2X1TS U2538 ( .A(n3272), .B(n3273), .Y(n3271) );
  NAND2X1TS U2539 ( .A(n3274), .B(n3275), .Y(n2968) );
  NAND2X1TS U2540 ( .A(n3278), .B(n3279), .Y(n3277) );
  NAND2X1TS U2541 ( .A(n2867), .B(n2798), .Y(n3279) );
  NAND2X1TS U2542 ( .A(n2846), .B(n2877), .Y(n3278) );
  NAND2X1TS U2543 ( .A(n3280), .B(n3281), .Y(n3276) );
  NAND2X1TS U2544 ( .A(n2764), .B(n2881), .Y(n3281) );
  NAND2X1TS U2545 ( .A(n3285), .B(n3286), .Y(n3284) );
  NAND2X1TS U2546 ( .A(n2848), .B(n3287), .Y(n3286) );
  NAND2X1TS U2547 ( .A(n3104), .B(n2739), .Y(n3287) );
  NAND2X1TS U2548 ( .A(n3161), .B(n3132), .Y(n3285) );
  NAND2X1TS U2549 ( .A(n3290), .B(n3291), .Y(n3283) );
  NAND2X1TS U2550 ( .A(n2841), .B(n3292), .Y(n3291) );
  NAND2X1TS U2551 ( .A(n2837), .B(n2823), .Y(n3292) );
  NAND2X1TS U2552 ( .A(n3296), .B(n3297), .Y(n2957) );
  NAND2X1TS U2553 ( .A(n3302), .B(n3303), .Y(n3301) );
  NAND2X1TS U2554 ( .A(n3304), .B(n2878), .Y(n3303) );
  NAND2X1TS U2555 ( .A(n2765), .B(n2986), .Y(n3302) );
  NAND2X1TS U2556 ( .A(n3307), .B(n3308), .Y(n3306) );
  NAND2X1TS U2557 ( .A(n3313), .B(n3314), .Y(n3305) );
  NAND2X1TS U2558 ( .A(n2781), .B(n2728), .Y(n3257) );
  NAND2X1TS U2559 ( .A(n2960), .B(n3323), .Y(n3322) );
  NAND2X1TS U2560 ( .A(n3328), .B(n3329), .Y(n3327) );
  NAND2X1TS U2561 ( .A(n2701), .B(n2737), .Y(n3329) );
  NAND2X1TS U2562 ( .A(n2854), .B(n3330), .Y(n3328) );
  NAND2X1TS U2563 ( .A(n3331), .B(n3332), .Y(n3326) );
  NAND2X1TS U2564 ( .A(n2858), .B(n3333), .Y(n3332) );
  NAND2X1TS U2565 ( .A(n2977), .B(n2830), .Y(n3333) );
  NAND2X1TS U2566 ( .A(n3338), .B(n3339), .Y(n3019) );
  NAND2X1TS U2567 ( .A(n3240), .B(n3342), .Y(n3341) );
  NAND2X1TS U2568 ( .A(n2886), .B(n2769), .Y(n3342) );
  NAND2X1TS U2569 ( .A(n3023), .B(n2786), .Y(n3240) );
  NAND2X1TS U2570 ( .A(n3343), .B(n3344), .Y(n3340) );
  NAND2X1TS U2571 ( .A(n3097), .B(n3330), .Y(n3344) );
  NAND2X1TS U2572 ( .A(n2704), .B(n2742), .Y(n3330) );
  NAND2X1TS U2573 ( .A(n2857), .B(n2763), .Y(n3343) );
  NAND2X1TS U2574 ( .A(n3347), .B(n3348), .Y(n3346) );
  NAND2X1TS U2575 ( .A(n2809), .B(n3349), .Y(n3348) );
  NAND2X1TS U2576 ( .A(n3350), .B(n2781), .Y(n3349) );
  NAND2X1TS U2577 ( .A(n2877), .B(n3351), .Y(n3347) );
  NAND2X1TS U2578 ( .A(n3169), .B(n2802), .Y(n3351) );
  NAND2X1TS U2579 ( .A(n3352), .B(n3353), .Y(n3345) );
  NAND2X1TS U2580 ( .A(n2924), .B(n3354), .Y(n3353) );
  NAND2X1TS U2581 ( .A(n2838), .B(n2767), .Y(n3354) );
  NAND2X1TS U2582 ( .A(n2744), .B(n3355), .Y(n3352) );
  NAND2X1TS U2583 ( .A(n3295), .B(n2831), .Y(n3355) );
  NAND2X1TS U2584 ( .A(n2707), .B(n3460), .Y(n3013) );
  NAND2X1TS U2585 ( .A(n2820), .B(n2792), .Y(n3356) );
  NAND2X1TS U2586 ( .A(n3359), .B(n3360), .Y(n3358) );
  NAND2X1TS U2587 ( .A(n2798), .B(n3361), .Y(n3360) );
  NAND2X1TS U2588 ( .A(n2800), .B(n2757), .Y(n3361) );
  NAND2X1TS U2589 ( .A(n2911), .B(n2908), .Y(n3573) );
  NAND2X1TS U2590 ( .A(n2726), .B(n3362), .Y(n3359) );
  NAND2X1TS U2591 ( .A(n2829), .B(n2735), .Y(n3362) );
  NAND2X1TS U2592 ( .A(n3366), .B(n3367), .Y(n3365) );
  NAND2X1TS U2593 ( .A(n2844), .B(n2865), .Y(n3367) );
  NAND2X1TS U2594 ( .A(n3370), .B(n2897), .Y(n3167) );
  NAND2X1TS U2595 ( .A(n3373), .B(n3374), .Y(n3372) );
  NAND2X1TS U2596 ( .A(n3499), .B(n2706), .Y(n2988) );
  NAND2X1TS U2597 ( .A(n3379), .B(n3244), .Y(n3378) );
  NAND2X1TS U2598 ( .A(n2869), .B(n2851), .Y(n3244) );
  NAND2X1TS U2599 ( .A(n2881), .B(n2848), .Y(n3379) );
  NAND2X1TS U2600 ( .A(n3459), .B(n2709), .Y(n3125) );
  NAND2X1TS U2601 ( .A(n3380), .B(n3381), .Y(n3371) );
  NAND2X1TS U2602 ( .A(n3387), .B(n3388), .Y(n3386) );
  NAND2X1TS U2603 ( .A(n2866), .B(n3389), .Y(n3388) );
  NAND2X1TS U2604 ( .A(n2794), .B(n2829), .Y(n3389) );
  NAND2X1TS U2605 ( .A(n3459), .B(n3428), .Y(n3089) );
  NAND2X1TS U2606 ( .A(n2874), .B(n3258), .Y(n3387) );
  NAND2X1TS U2607 ( .A(n2795), .B(n2723), .Y(n3258) );
  NAND2X1TS U2608 ( .A(n2740), .B(n2838), .Y(n3115) );
  NAND2X1TS U2609 ( .A(n2730), .B(n2845), .Y(n3391) );
  NAND2X1TS U2610 ( .A(n3394), .B(n3395), .Y(n3393) );
  NAND2X1TS U2611 ( .A(n2714), .B(n3396), .Y(n3395) );
  NAND2X1TS U2612 ( .A(n2837), .B(n2715), .Y(n3396) );
  NAND2X1TS U2613 ( .A(n3560), .B(n3561), .Y(n2954) );
  NAND2X1TS U2614 ( .A(n2698), .B(n3397), .Y(n3394) );
  NAND2X1TS U2615 ( .A(n3398), .B(n2772), .Y(n3397) );
  NAND2X1TS U2616 ( .A(n3399), .B(n3400), .Y(n3392) );
  NAND2X1TS U2617 ( .A(n2725), .B(n3401), .Y(n3400) );
  NAND2X1TS U2618 ( .A(n2793), .B(n2806), .Y(n3401) );
  NAND2X1TS U2619 ( .A(n3408), .B(n3409), .Y(n3407) );
  NAND2X1TS U2620 ( .A(n2707), .B(n3428), .Y(n3096) );
  NAND2X1TS U2621 ( .A(n3414), .B(n3415), .Y(n3406) );
  NAND2X1TS U2622 ( .A(n2697), .B(n2722), .Y(n3288) );
  NAND2X1TS U2623 ( .A(n2899), .B(n3586), .Y(n3398) );
  NAND2X1TS U2624 ( .A(n2912), .B(n2895), .Y(n3527) );
  NAND2X1TS U2625 ( .A(n3422), .B(n3423), .Y(n3421) );
  NAND2X1TS U2626 ( .A(n2738), .B(n3424), .Y(n3423) );
  NAND2X1TS U2627 ( .A(n2801), .B(n2719), .Y(n3424) );
  NAND2X1TS U2628 ( .A(n2909), .B(n2889), .Y(n3524) );
  NAND2X1TS U2629 ( .A(n3555), .B(n3459), .Y(n3080) );
  NAND2X1TS U2630 ( .A(n2854), .B(n3425), .Y(n3422) );
  NAND2X1TS U2631 ( .A(n2801), .B(n2780), .Y(n3425) );
  NAND2X1TS U2632 ( .A(n2911), .B(n3570), .Y(n3569) );
  NAND2X1TS U2633 ( .A(n2893), .B(n3428), .Y(n3427) );
  MXI2X1TS U2634 ( .A(n3429), .B(n2744), .S0(n2905), .Y(n3426) );
  NAND2X1TS U2635 ( .A(n3560), .B(n3587), .Y(n2945) );
  NAND2X1TS U2636 ( .A(n2728), .B(n2824), .Y(n3429) );
  NAND2X1TS U2637 ( .A(n2895), .B(n3562), .Y(n3578) );
endmodule

