%%% protect protected_file
module AND2 (
  Y,
  A,
  B
)
;
output Y ;
input A ;
input B ;
endmodule /* AND2 */

module AND2A (
  Y,
  A,
  B
)
;
output Y ;
input A ;
input B ;
endmodule /* AND2A */

module AND2B (
  Y,
  A,
  B
)
;
output Y ;
input A ;
input B ;
endmodule /* AND2B */

module AND3 (
  Y,
  A,
  B,
  C
)
;
output Y ;
input A ;
input B ;
input C ;
endmodule /* AND3 */

module AND3A (
  Y,
  A,
  B,
  C
)
;
output Y ;
input A ;
input B ;
input C ;
endmodule /* AND3A */

module AND3B (
  Y,
  A,
  B,
  C
)
;
output Y ;
input A ;
input B ;
input C ;
endmodule /* AND3B */

module AND3C (
  Y,
  A,
  B,
  C
)
;
output Y ;
input A ;
input B ;
input C ;
endmodule /* AND3C */

module AO1 (
  Y,
  A,
  B,
  C
)
;
output Y ;
input A ;
input B ;
input C ;
endmodule /* AO1 */

module AO12 (
  Y,
  A,
  B,
  C
)
;
output Y ;
input A ;
input B ;
input C ;
endmodule /* AO12 */

module AO13 (
  Y,
  A,
  B,
  C
)
;
output Y ;
input A ;
input B ;
input C ;
endmodule /* AO13 */

module AO14 (
  Y,
  A,
  B,
  C
)
;
output Y ;
input A ;
input B ;
input C ;
endmodule /* AO14 */

module AO15 (
  Y,
  A,
  B,
  C
)
;
output Y ;
input A ;
input B ;
input C ;
endmodule /* AO15 */

module AO16 (
  Y,
  A,
  B,
  C
)
;
output Y ;
input A ;
input B ;
input C ;
endmodule /* AO16 */

module AO17 (
  Y,
  A,
  B,
  C
)
;
output Y ;
input A ;
input B ;
input C ;
endmodule /* AO17 */

module AO18 (
  Y,
  A,
  B,
  C
)
;
output Y ;
input A ;
input B ;
input C ;
endmodule /* AO18 */

module AO1A (
  Y,
  A,
  B,
  C
)
;
output Y ;
input A ;
input B ;
input C ;
endmodule /* AO1A */

module AO1B (
  Y,
  A,
  B,
  C
)
;
output Y ;
input A ;
input B ;
input C ;
endmodule /* AO1B */

module AO1C (
  Y,
  A,
  B,
  C
)
;
output Y ;
input A ;
input B ;
input C ;
endmodule /* AO1C */

module AO1D (
  Y,
  A,
  B,
  C
)
;
output Y ;
input A ;
input B ;
input C ;
endmodule /* AO1D */

module AO1E (
  Y,
  A,
  B,
  C
)
;
output Y ;
input A ;
input B ;
input C ;
endmodule /* AO1E */

module AOI1 (
  Y,
  A,
  B,
  C
)
;
output Y ;
input A ;
input B ;
input C ;
endmodule /* AOI1 */

module AOI1A (
  Y,
  A,
  B,
  C
)
;
output Y ;
input A ;
input B ;
input C ;
endmodule /* AOI1A */

module AOI1B (
  Y,
  A,
  B,
  C
)
;
output Y ;
input A ;
input B ;
input C ;
endmodule /* AOI1B */

module AOI1C (
  Y,
  A,
  B,
  C
)
;
output Y ;
input A ;
input B ;
input C ;
endmodule /* AOI1C */

module AOI1D (
  Y,
  A,
  B,
  C
)
;
output Y ;
input A ;
input B ;
input C ;
endmodule /* AOI1D */

module AOI5 (
  Y,
  A,
  B,
  C
)
;
output Y ;
input A ;
input B ;
input C ;
endmodule /* AOI5 */

module AX1 (
  Y,
  A,
  B,
  C
)
;
output Y ;
input A ;
input B ;
input C ;
endmodule /* AX1 */

module AX1A (
  Y,
  A,
  B,
  C
)
;
output Y ;
input A ;
input B ;
input C ;
endmodule /* AX1A */

module AX1B (
  Y,
  A,
  B,
  C
)
;
output Y ;
input A ;
input B ;
input C ;
endmodule /* AX1B */

module AX1C (
  Y,
  A,
  B,
  C
)
;
output Y ;
input A ;
input B ;
input C ;
endmodule /* AX1C */

module AX1D (
  Y,
  A,
  B,
  C
)
;
output Y ;
input A ;
input B ;
input C ;
endmodule /* AX1D */

module AX1E (
  Y,
  A,
  B,
  C
)
;
output Y ;
input A ;
input B ;
input C ;
endmodule /* AX1E */

module AXO1 (
  Y,
  A,
  B,
  C
)
;
output Y ;
input A ;
input B ;
input C ;
endmodule /* AXO1 */

module AXO2 (
  Y,
  A,
  B,
  C
)
;
output Y ;
input A ;
input B ;
input C ;
endmodule /* AXO2 */

module AXO3 (
  Y,
  A,
  B,
  C
)
;
output Y ;
input A ;
input B ;
input C ;
endmodule /* AXO3 */

module AXO5 (
  Y,
  A,
  B,
  C
)
;
output Y ;
input A ;
input B ;
input C ;
endmodule /* AXO5 */

module AXO6 (
  Y,
  A,
  B,
  C
)
;
output Y ;
input A ;
input B ;
input C ;
endmodule /* AXO6 */

module AXO7 (
  Y,
  A,
  B,
  C
)
;
output Y ;
input A ;
input B ;
input C ;
endmodule /* AXO7 */

module AXOI1 (
  Y,
  A,
  B,
  C
)
;
output Y ;
input A ;
input B ;
input C ;
endmodule /* AXOI1 */

module AXOI2 (
  Y,
  A,
  B,
  C
)
;
output Y ;
input A ;
input B ;
input C ;
endmodule /* AXOI2 */

module AXOI3 (
  Y,
  A,
  B,
  C
)
;
output Y ;
input A ;
input B ;
input C ;
endmodule /* AXOI3 */

module AXOI4 (
  Y,
  A,
  B,
  C
)
;
output Y ;
input A ;
input B ;
input C ;
endmodule /* AXOI4 */

module AXOI5 (
  Y,
  A,
  B,
  C
)
;
output Y ;
input A ;
input B ;
input C ;
endmodule /* AXOI5 */

module AXOI7 (
  Y,
  A,
  B,
  C
)
;
output Y ;
input A ;
input B ;
input C ;
endmodule /* AXOI7 */

module BIBUF (
  PAD,
  Y,
  D,
  E
)
;
inout PAD /* synthesis syn_tristate = 1 */ ;
output Y ;
input D ;
input E ;
endmodule /* BIBUF */

module BIBUF_F_2 (
  PAD,
  Y,
  D,
  E
)
;
inout PAD /* synthesis syn_tristate = 1 */ ;
output Y ;
input D ;
input E ;
endmodule /* BIBUF_F_2 */

module BIBUF_F_2D (
  PAD,
  Y,
  D,
  E
)
;
inout PAD /* synthesis syn_tristate = 1 */ ;
output Y ;
input D ;
input E ;
endmodule /* BIBUF_F_2D */

module BIBUF_F_2U (
  PAD,
  Y,
  D,
  E
)
;
inout PAD /* synthesis syn_tristate = 1 */ ;
output Y ;
input D ;
input E ;
endmodule /* BIBUF_F_2U */

module BIBUF_F_4 (
  PAD,
  Y,
  D,
  E
)
;
inout PAD /* synthesis syn_tristate = 1 */ ;
output Y ;
input D ;
input E ;
endmodule /* BIBUF_F_4 */

module BIBUF_F_4D (
  PAD,
  Y,
  D,
  E
)
;
inout PAD /* synthesis syn_tristate = 1 */ ;
output Y ;
input D ;
input E ;
endmodule /* BIBUF_F_4D */

module BIBUF_F_4U (
  PAD,
  Y,
  D,
  E
)
;
inout PAD /* synthesis syn_tristate = 1 */ ;
output Y ;
input D ;
input E ;
endmodule /* BIBUF_F_4U */

module BIBUF_F_6 (
  PAD,
  Y,
  D,
  E
)
;
inout PAD /* synthesis syn_tristate = 1 */ ;
output Y ;
input D ;
input E ;
endmodule /* BIBUF_F_6 */

module BIBUF_F_6D (
  PAD,
  Y,
  D,
  E
)
;
inout PAD /* synthesis syn_tristate = 1 */ ;
output Y ;
input D ;
input E ;
endmodule /* BIBUF_F_6D */

module BIBUF_F_6U (
  PAD,
  Y,
  D,
  E
)
;
inout PAD /* synthesis syn_tristate = 1 */ ;
output Y ;
input D ;
input E ;
endmodule /* BIBUF_F_6U */

module BIBUF_F_8 (
  PAD,
  Y,
  D,
  E
)
;
inout PAD /* synthesis syn_tristate = 1 */ ;
output Y ;
input D ;
input E ;
endmodule /* BIBUF_F_8 */

module BIBUF_F_8D (
  PAD,
  Y,
  D,
  E
)
;
inout PAD /* synthesis syn_tristate = 1 */ ;
output Y ;
input D ;
input E ;
endmodule /* BIBUF_F_8D */

module BIBUF_F_8U (
  PAD,
  Y,
  D,
  E
)
;
inout PAD /* synthesis syn_tristate = 1 */ ;
output Y ;
input D ;
input E ;
endmodule /* BIBUF_F_8U */

module BIBUF_F_12 (
  PAD,
  Y,
  D,
  E
)
;
inout PAD /* synthesis syn_tristate = 1 */ ;
output Y ;
input D ;
input E ;
endmodule /* BIBUF_F_12 */

module BIBUF_F_12D (
  PAD,
  Y,
  D,
  E
)
;
inout PAD /* synthesis syn_tristate = 1 */ ;
output Y ;
input D ;
input E ;
endmodule /* BIBUF_F_12D */

module BIBUF_F_12U (
  PAD,
  Y,
  D,
  E
)
;
inout PAD /* synthesis syn_tristate = 1 */ ;
output Y ;
input D ;
input E ;
endmodule /* BIBUF_F_12U */

module BIBUF_F_16 (
  PAD,
  Y,
  D,
  E
)
;
inout PAD /* synthesis syn_tristate = 1 */ ;
output Y ;
input D ;
input E ;
endmodule /* BIBUF_F_16 */

module BIBUF_F_16D (
  PAD,
  Y,
  D,
  E
)
;
inout PAD /* synthesis syn_tristate = 1 */ ;
output Y ;
input D ;
input E ;
endmodule /* BIBUF_F_16D */

module BIBUF_F_16U (
  PAD,
  Y,
  D,
  E
)
;
inout PAD /* synthesis syn_tristate = 1 */ ;
output Y ;
input D ;
input E ;
endmodule /* BIBUF_F_16U */

module BIBUF_F_24 (
  PAD,
  Y,
  D,
  E
)
;
inout PAD /* synthesis syn_tristate = 1 */ ;
output Y ;
input D ;
input E ;
endmodule /* BIBUF_F_24 */

module BIBUF_F_24D (
  PAD,
  Y,
  D,
  E
)
;
inout PAD /* synthesis syn_tristate = 1 */ ;
output Y ;
input D ;
input E ;
endmodule /* BIBUF_F_24D */

module BIBUF_F_24U (
  PAD,
  Y,
  D,
  E
)
;
inout PAD /* synthesis syn_tristate = 1 */ ;
output Y ;
input D ;
input E ;
endmodule /* BIBUF_F_24U */

module BIBUF_GTL25 (
  PAD,
  Y,
  D,
  E
)
;
inout PAD /* synthesis syn_tristate = 1 */ ;
output Y ;
input D ;
input E ;
endmodule /* BIBUF_GTL25 */

module BIBUF_GTL33 (
  PAD,
  Y,
  D,
  E
)
;
inout PAD /* synthesis syn_tristate = 1 */ ;
output Y ;
input D ;
input E ;
endmodule /* BIBUF_GTL33 */

module BIBUF_GTLP25 (
  PAD,
  Y,
  D,
  E
)
;
inout PAD /* synthesis syn_tristate = 1 */ ;
output Y ;
input D ;
input E ;
endmodule /* BIBUF_GTLP25 */

module BIBUF_GTLP33 (
  PAD,
  Y,
  D,
  E
)
;
inout PAD /* synthesis syn_tristate = 1 */ ;
output Y ;
input D ;
input E ;
endmodule /* BIBUF_GTLP33 */

module BIBUF_HSTL_I (
  PAD,
  Y,
  D,
  E
)
;
inout PAD /* synthesis syn_tristate = 1 */ ;
output Y ;
input D ;
input E ;
endmodule /* BIBUF_HSTL_I */

module BIBUF_HSTL_II (
  PAD,
  Y,
  D,
  E
)
;
inout PAD /* synthesis syn_tristate = 1 */ ;
output Y ;
input D ;
input E ;
endmodule /* BIBUF_HSTL_II */

module BIBUF_LVCMOS15 (
  PAD,
  Y,
  D,
  E
)
;
inout PAD /* synthesis syn_tristate = 1 */ ;
output Y ;
input D ;
input E ;
endmodule /* BIBUF_LVCMOS15 */

module BIBUF_LVCMOS15D (
  PAD,
  Y,
  D,
  E
)
;
inout PAD /* synthesis syn_tristate = 1 */ ;
output Y ;
input D ;
input E ;
endmodule /* BIBUF_LVCMOS15D */

module BIBUF_LVCMOS15U (
  PAD,
  Y,
  D,
  E
)
;
inout PAD /* synthesis syn_tristate = 1 */ ;
output Y ;
input D ;
input E ;
endmodule /* BIBUF_LVCMOS15U */

module BIBUF_LVCMOS18 (
  PAD,
  Y,
  D,
  E
)
;
inout PAD /* synthesis syn_tristate = 1 */ ;
output Y ;
input D ;
input E ;
endmodule /* BIBUF_LVCMOS18 */

module BIBUF_LVCMOS18D (
  PAD,
  Y,
  D,
  E
)
;
inout PAD /* synthesis syn_tristate = 1 */ ;
output Y ;
input D ;
input E ;
endmodule /* BIBUF_LVCMOS18D */

module BIBUF_LVCMOS18U (
  PAD,
  Y,
  D,
  E
)
;
inout PAD /* synthesis syn_tristate = 1 */ ;
output Y ;
input D ;
input E ;
endmodule /* BIBUF_LVCMOS18U */

module BIBUF_LVCMOS25 (
  PAD,
  Y,
  D,
  E
)
;
inout PAD /* synthesis syn_tristate = 1 */ ;
output Y ;
input D ;
input E ;
endmodule /* BIBUF_LVCMOS25 */

module BIBUF_LVCMOS25D (
  PAD,
  Y,
  D,
  E
)
;
inout PAD /* synthesis syn_tristate = 1 */ ;
output Y ;
input D ;
input E ;
endmodule /* BIBUF_LVCMOS25D */

module BIBUF_LVCMOS25U (
  PAD,
  Y,
  D,
  E
)
;
inout PAD /* synthesis syn_tristate = 1 */ ;
output Y ;
input D ;
input E ;
endmodule /* BIBUF_LVCMOS25U */

module BIBUF_LVCMOS33 (
  PAD,
  Y,
  D,
  E
)
;
inout PAD /* synthesis syn_tristate = 1 */ ;
output Y ;
input D ;
input E ;
endmodule /* BIBUF_LVCMOS33 */

module BIBUF_LVCMOS33D (
  PAD,
  Y,
  D,
  E
)
;
inout PAD /* synthesis syn_tristate = 1 */ ;
output Y ;
input D ;
input E ;
endmodule /* BIBUF_LVCMOS33D */

module BIBUF_LVCMOS33U (
  PAD,
  Y,
  D,
  E
)
;
inout PAD /* synthesis syn_tristate = 1 */ ;
output Y ;
input D ;
input E ;
endmodule /* BIBUF_LVCMOS33U */

module BIBUF_LVCMOS5 (
  PAD,
  Y,
  D,
  E
)
;
inout PAD /* synthesis syn_tristate = 1 */ ;
output Y ;
input D ;
input E ;
endmodule /* BIBUF_LVCMOS5 */

module BIBUF_LVCMOS5D (
  PAD,
  Y,
  D,
  E
)
;
inout PAD /* synthesis syn_tristate = 1 */ ;
output Y ;
input D ;
input E ;
endmodule /* BIBUF_LVCMOS5D */

module BIBUF_LVCMOS5U (
  PAD,
  Y,
  D,
  E
)
;
inout PAD /* synthesis syn_tristate = 1 */ ;
output Y ;
input D ;
input E ;
endmodule /* BIBUF_LVCMOS5U */

module BIBUF_PCI (
  PAD,
  Y,
  D,
  E
)
;
inout PAD /* synthesis syn_tristate = 1 */ ;
output Y ;
input D ;
input E ;
endmodule /* BIBUF_PCI */

module BIBUF_PCIX (
  PAD,
  Y,
  D,
  E
)
;
inout PAD /* synthesis syn_tristate = 1 */ ;
output Y ;
input D ;
input E ;
endmodule /* BIBUF_PCIX */

module BIBUF_S_2 (
  PAD,
  Y,
  D,
  E
)
;
inout PAD /* synthesis syn_tristate = 1 */ ;
output Y ;
input D ;
input E ;
endmodule /* BIBUF_S_2 */

module BIBUF_S_2D (
  PAD,
  Y,
  D,
  E
)
;
inout PAD /* synthesis syn_tristate = 1 */ ;
output Y ;
input D ;
input E ;
endmodule /* BIBUF_S_2D */

module BIBUF_S_2U (
  PAD,
  Y,
  D,
  E
)
;
inout PAD /* synthesis syn_tristate = 1 */ ;
output Y ;
input D ;
input E ;
endmodule /* BIBUF_S_2U */

module BIBUF_S_4 (
  PAD,
  Y,
  D,
  E
)
;
inout PAD /* synthesis syn_tristate = 1 */ ;
output Y ;
input D ;
input E ;
endmodule /* BIBUF_S_4 */

module BIBUF_S_4D (
  PAD,
  Y,
  D,
  E
)
;
inout PAD /* synthesis syn_tristate = 1 */ ;
output Y ;
input D ;
input E ;
endmodule /* BIBUF_S_4D */

module BIBUF_S_4U (
  PAD,
  Y,
  D,
  E
)
;
inout PAD /* synthesis syn_tristate = 1 */ ;
output Y ;
input D ;
input E ;
endmodule /* BIBUF_S_4U */

module BIBUF_S_6 (
  PAD,
  Y,
  D,
  E
)
;
inout PAD /* synthesis syn_tristate = 1 */ ;
output Y ;
input D ;
input E ;
endmodule /* BIBUF_S_6 */

module BIBUF_S_6D (
  PAD,
  Y,
  D,
  E
)
;
inout PAD /* synthesis syn_tristate = 1 */ ;
output Y ;
input D ;
input E ;
endmodule /* BIBUF_S_6D */

module BIBUF_S_6U (
  PAD,
  Y,
  D,
  E
)
;
inout PAD /* synthesis syn_tristate = 1 */ ;
output Y ;
input D ;
input E ;
endmodule /* BIBUF_S_6U */

module BIBUF_S_8 (
  PAD,
  Y,
  D,
  E
)
;
inout PAD /* synthesis syn_tristate = 1 */ ;
output Y ;
input D ;
input E ;
endmodule /* BIBUF_S_8 */

module BIBUF_S_8D (
  PAD,
  Y,
  D,
  E
)
;
inout PAD /* synthesis syn_tristate = 1 */ ;
output Y ;
input D ;
input E ;
endmodule /* BIBUF_S_8D */

module BIBUF_S_8U (
  PAD,
  Y,
  D,
  E
)
;
inout PAD /* synthesis syn_tristate = 1 */ ;
output Y ;
input D ;
input E ;
endmodule /* BIBUF_S_8U */

module BIBUF_S_12 (
  PAD,
  Y,
  D,
  E
)
;
inout PAD /* synthesis syn_tristate = 1 */ ;
output Y ;
input D ;
input E ;
endmodule /* BIBUF_S_12 */

module BIBUF_S_12D (
  PAD,
  Y,
  D,
  E
)
;
inout PAD /* synthesis syn_tristate = 1 */ ;
output Y ;
input D ;
input E ;
endmodule /* BIBUF_S_12D */

module BIBUF_S_12U (
  PAD,
  Y,
  D,
  E
)
;
inout PAD /* synthesis syn_tristate = 1 */ ;
output Y ;
input D ;
input E ;
endmodule /* BIBUF_S_12U */

module BIBUF_S_16 (
  PAD,
  Y,
  D,
  E
)
;
inout PAD /* synthesis syn_tristate = 1 */ ;
output Y ;
input D ;
input E ;
endmodule /* BIBUF_S_16 */

module BIBUF_S_16D (
  PAD,
  Y,
  D,
  E
)
;
inout PAD /* synthesis syn_tristate = 1 */ ;
output Y ;
input D ;
input E ;
endmodule /* BIBUF_S_16D */

module BIBUF_S_16U (
  PAD,
  Y,
  D,
  E
)
;
inout PAD /* synthesis syn_tristate = 1 */ ;
output Y ;
input D ;
input E ;
endmodule /* BIBUF_S_16U */

module BIBUF_S_24 (
  PAD,
  Y,
  D,
  E
)
;
inout PAD /* synthesis syn_tristate = 1 */ ;
output Y ;
input D ;
input E ;
endmodule /* BIBUF_S_24 */

module BIBUF_S_24D (
  PAD,
  Y,
  D,
  E
)
;
inout PAD /* synthesis syn_tristate = 1 */ ;
output Y ;
input D ;
input E ;
endmodule /* BIBUF_S_24D */

module BIBUF_S_24U (
  PAD,
  Y,
  D,
  E
)
;
inout PAD /* synthesis syn_tristate = 1 */ ;
output Y ;
input D ;
input E ;
endmodule /* BIBUF_S_24U */

module BIBUF_SSTL2_I (
  PAD,
  Y,
  D,
  E
)
;
inout PAD /* synthesis syn_tristate = 1 */ ;
output Y ;
input D ;
input E ;
endmodule /* BIBUF_SSTL2_I */

module BIBUF_SSTL2_II (
  PAD,
  Y,
  D,
  E
)
;
inout PAD /* synthesis syn_tristate = 1 */ ;
output Y ;
input D ;
input E ;
endmodule /* BIBUF_SSTL2_II */

module BIBUF_SSTL3_I (
  PAD,
  Y,
  D,
  E
)
;
inout PAD /* synthesis syn_tristate = 1 */ ;
output Y ;
input D ;
input E ;
endmodule /* BIBUF_SSTL3_I */

module BIBUF_SSTL3_II (
  PAD,
  Y,
  D,
  E
)
;
inout PAD /* synthesis syn_tristate = 1 */ ;
output Y ;
input D ;
input E ;
endmodule /* BIBUF_SSTL3_II */

module BIBUF_LVDS (
  PADN,
  PADP,
  Y,
  D,
  E
)
;
inout PADN /* synthesis syn_tristate = 1 */ ;
inout PADP /* synthesis syn_tristate = 1 */ ;
output Y ;
input D ;
input E ;
endmodule /* BIBUF_LVDS */

module BUFD (
  Y,
  A
)
;
output Y ;
input A ;
endmodule /* BUFD */

module BUFF (
  Y,
  A
)
;
output Y ;
input A ;
endmodule /* BUFF */

module CLKBIBUF (
  PAD,
  Y,
  D,
  E
)
;
inout PAD /* synthesis syn_tristate = 1 */ ;
output Y ;
input D ;
input E ;
endmodule /* CLKBIBUF */

module CLKBUF (
  Y,
  PAD
)
;
output Y ;
input PAD ;
endmodule /* CLKBUF */

module CLKBUF_GTL25 (
  Y,
  PAD
)
;
output Y ;
input PAD ;
endmodule /* CLKBUF_GTL25 */

module CLKBUF_GTL33 (
  Y,
  PAD
)
;
output Y ;
input PAD ;
endmodule /* CLKBUF_GTL33 */

module CLKBUF_GTLP25 (
  Y,
  PAD
)
;
output Y ;
input PAD ;
endmodule /* CLKBUF_GTLP25 */

module CLKBUF_GTLP33 (
  Y,
  PAD
)
;
output Y ;
input PAD ;
endmodule /* CLKBUF_GTLP33 */

module CLKBUF_HSTL_I (
  Y,
  PAD
)
;
output Y ;
input PAD ;
endmodule /* CLKBUF_HSTL_I */

module CLKBUF_HSTL_II (
  Y,
  PAD
)
;
output Y ;
input PAD ;
endmodule /* CLKBUF_HSTL_II */

module CLKBUF_LVCMOS15 (
  Y,
  PAD
)
;
output Y ;
input PAD ;
endmodule /* CLKBUF_LVCMOS15 */

module CLKBUF_LVCMOS18 (
  Y,
  PAD
)
;
output Y ;
input PAD ;
endmodule /* CLKBUF_LVCMOS18 */

module CLKBUF_LVCMOS25 (
  Y,
  PAD
)
;
output Y ;
input PAD ;
endmodule /* CLKBUF_LVCMOS25 */

module CLKBUF_LVCMOS33 (
  Y,
  PAD
)
;
output Y ;
input PAD ;
endmodule /* CLKBUF_LVCMOS33 */

module CLKBUF_LVCMOS5 (
  Y,
  PAD
)
;
output Y ;
input PAD ;
endmodule /* CLKBUF_LVCMOS5 */

module CLKBUF_PCI (
  Y,
  PAD
)
;
output Y ;
input PAD ;
endmodule /* CLKBUF_PCI */

module CLKBUF_PCIX (
  Y,
  PAD
)
;
output Y ;
input PAD ;
endmodule /* CLKBUF_PCIX */

module CLKBUF_SSTL2_I (
  Y,
  PAD
)
;
output Y ;
input PAD ;
endmodule /* CLKBUF_SSTL2_I */

module CLKBUF_SSTL2_II (
  Y,
  PAD
)
;
output Y ;
input PAD ;
endmodule /* CLKBUF_SSTL2_II */

module CLKBUF_SSTL3_I (
  Y,
  PAD
)
;
output Y ;
input PAD ;
endmodule /* CLKBUF_SSTL3_I */

module CLKBUF_SSTL3_II (
  Y,
  PAD
)
;
output Y ;
input PAD ;
endmodule /* CLKBUF_SSTL3_II */

module CLKINT (
  Y,
  A
)
;
output Y ;
input A ;
endmodule /* CLKINT */

module CLKIO (
  Y,
  A
)
;
output Y ;
input A ;
endmodule /* CLKIO */

module DFI0 (
  QN,
  CLK,
  D
)
;
output QN ;
input CLK ;
input D ;
endmodule /* DFI0 */

module DFI0C0 (
  QN,
  CLK,
  CLR,
  D
)
;
output QN ;
input CLK ;
input CLR ;
input D ;
endmodule /* DFI0C0 */

module DFI0C1 (
  QN,
  CLK,
  CLR,
  D
)
;
output QN ;
input CLK ;
input CLR ;
input D ;
endmodule /* DFI0C1 */

module DFI0E0 (
  QN,
  CLK,
  D,
  E
)
;
output QN ;
input CLK ;
input D ;
input E ;
endmodule /* DFI0E0 */

module DFI0E0C0 (
  QN,
  CLK,
  CLR,
  D,
  E
)
;
output QN ;
input CLK ;
input CLR ;
input D ;
input E ;
endmodule /* DFI0E0C0 */

module DFI0E0C1 (
  QN,
  CLK,
  CLR,
  D,
  E
)
;
output QN ;
input CLK ;
input CLR ;
input D ;
input E ;
endmodule /* DFI0E0C1 */

module DFI0E0P0 (
  QN,
  CLK,
  D,
  E,
  PRE
)
;
output QN ;
input CLK ;
input D ;
input E ;
input PRE ;
endmodule /* DFI0E0P0 */

module DFI0E0P1 (
  QN,
  CLK,
  D,
  E,
  PRE
)
;
output QN ;
input CLK ;
input D ;
input E ;
input PRE ;
endmodule /* DFI0E0P1 */

module DFI0E1 (
  QN,
  CLK,
  D,
  E
)
;
output QN ;
input CLK ;
input D ;
input E ;
endmodule /* DFI0E1 */

module DFI0E1C0 (
  QN,
  CLK,
  CLR,
  D,
  E
)
;
output QN ;
input CLK ;
input CLR ;
input D ;
input E ;
endmodule /* DFI0E1C0 */

module DFI0E1C1 (
  QN,
  CLK,
  CLR,
  D,
  E
)
;
output QN ;
input CLK ;
input CLR ;
input D ;
input E ;
endmodule /* DFI0E1C1 */

module DFI0E1P0 (
  QN,
  CLK,
  D,
  E,
  PRE
)
;
output QN ;
input CLK ;
input D ;
input E ;
input PRE ;
endmodule /* DFI0E1P0 */

module DFI0E1P1 (
  QN,
  CLK,
  D,
  E,
  PRE
)
;
output QN ;
input CLK ;
input D ;
input E ;
input PRE ;
endmodule /* DFI0E1P1 */

module DFI0P0 (
  QN,
  CLK,
  D,
  PRE
)
;
output QN ;
input CLK ;
input D ;
input PRE ;
endmodule /* DFI0P0 */

module DFI0P1 (
  QN,
  CLK,
  D,
  PRE
)
;
output QN ;
input CLK ;
input D ;
input PRE ;
endmodule /* DFI0P1 */

module DFI0P1C1 (
  QN,
  CLK,
  CLR,
  D,
  PRE
)
;
output QN ;
input CLK ;
input CLR ;
input D ;
input PRE ;
endmodule /* DFI0P1C1 */

module DFI1 (
  QN,
  CLK,
  D
)
;
output QN ;
input CLK ;
input D ;
endmodule /* DFI1 */

module DFI1C0 (
  QN,
  CLK,
  CLR,
  D
)
;
output QN ;
input CLK ;
input CLR ;
input D ;
endmodule /* DFI1C0 */

module DFI1C1 (
  QN,
  CLK,
  CLR,
  D
)
;
output QN ;
input CLK ;
input CLR ;
input D ;
endmodule /* DFI1C1 */

module DFI1E0 (
  QN,
  CLK,
  D,
  E
)
;
output QN ;
input CLK ;
input D ;
input E ;
endmodule /* DFI1E0 */

module DFI1E0C0 (
  QN,
  CLK,
  CLR,
  D,
  E
)
;
output QN ;
input CLK ;
input CLR ;
input D ;
input E ;
endmodule /* DFI1E0C0 */

module DFI1E0C1 (
  QN,
  CLK,
  CLR,
  D,
  E
)
;
output QN ;
input CLK ;
input CLR ;
input D ;
input E ;
endmodule /* DFI1E0C1 */

module DFI1E0P0 (
  QN,
  CLK,
  D,
  E,
  PRE
)
;
output QN ;
input CLK ;
input D ;
input E ;
input PRE ;
endmodule /* DFI1E0P0 */

module DFI1E0P1 (
  QN,
  CLK,
  D,
  E,
  PRE
)
;
output QN ;
input CLK ;
input D ;
input E ;
input PRE ;
endmodule /* DFI1E0P1 */

module DFI1E1 (
  QN,
  CLK,
  D,
  E
)
;
output QN ;
input CLK ;
input D ;
input E ;
endmodule /* DFI1E1 */

module DFI1E1C0 (
  QN,
  CLK,
  CLR,
  D,
  E
)
;
output QN ;
input CLK ;
input CLR ;
input D ;
input E ;
endmodule /* DFI1E1C0 */

module DFI1E1C1 (
  QN,
  CLK,
  CLR,
  D,
  E
)
;
output QN ;
input CLK ;
input CLR ;
input D ;
input E ;
endmodule /* DFI1E1C1 */

module DFI1E1P0 (
  QN,
  CLK,
  D,
  E,
  PRE
)
;
output QN ;
input CLK ;
input D ;
input E ;
input PRE ;
endmodule /* DFI1E1P0 */

module DFI1E1P1 (
  QN,
  CLK,
  D,
  E,
  PRE
)
;
output QN ;
input CLK ;
input D ;
input E ;
input PRE ;
endmodule /* DFI1E1P1 */

module DFI1P0 (
  QN,
  CLK,
  D,
  PRE
)
;
output QN ;
input CLK ;
input D ;
input PRE ;
endmodule /* DFI1P0 */

module DFI1P1 (
  QN,
  CLK,
  D,
  PRE
)
;
output QN ;
input CLK ;
input D ;
input PRE ;
endmodule /* DFI1P1 */

module DFI1P1C1 (
  QN,
  CLK,
  CLR,
  D,
  PRE
)
;
output QN ;
input CLK ;
input CLR ;
input D ;
input PRE ;
endmodule /* DFI1P1C1 */

module DFN0 (
  Q,
  CLK,
  D
)
;
output Q ;
input CLK ;
input D ;
endmodule /* DFN0 */

module DFN0C0 (
  Q,
  CLK,
  CLR,
  D
)
;
output Q ;
input CLK ;
input CLR ;
input D ;
endmodule /* DFN0C0 */

module DFN0C1 (
  Q,
  CLK,
  CLR,
  D
)
;
output Q ;
input CLK ;
input CLR ;
input D ;
endmodule /* DFN0C1 */

module DFN0E0 (
  Q,
  CLK,
  D,
  E
)
;
output Q ;
input CLK ;
input D ;
input E ;
endmodule /* DFN0E0 */

module DFN0E0C0 (
  Q,
  CLK,
  CLR,
  D,
  E
)
;
output Q ;
input CLK ;
input CLR ;
input D ;
input E ;
endmodule /* DFN0E0C0 */

module DFN0E0C1 (
  Q,
  CLK,
  CLR,
  D,
  E
)
;
output Q ;
input CLK ;
input CLR ;
input D ;
input E ;
endmodule /* DFN0E0C1 */

module DFN0E0P0 (
  Q,
  CLK,
  D,
  E,
  PRE
)
;
output Q ;
input CLK ;
input D ;
input E ;
input PRE ;
endmodule /* DFN0E0P0 */

module DFN0E0P1 (
  Q,
  CLK,
  D,
  E,
  PRE
)
;
output Q ;
input CLK ;
input D ;
input E ;
input PRE ;
endmodule /* DFN0E0P1 */

module DFN0E1 (
  Q,
  CLK,
  D,
  E
)
;
output Q ;
input CLK ;
input D ;
input E ;
endmodule /* DFN0E1 */

module DFN0E1C0 (
  Q,
  CLK,
  CLR,
  D,
  E
)
;
output Q ;
input CLK ;
input CLR ;
input D ;
input E ;
endmodule /* DFN0E1C0 */

module DFN0E1C1 (
  Q,
  CLK,
  CLR,
  D,
  E
)
;
output Q ;
input CLK ;
input CLR ;
input D ;
input E ;
endmodule /* DFN0E1C1 */

module DFN0E1P0 (
  Q,
  CLK,
  D,
  E,
  PRE
)
;
output Q ;
input CLK ;
input D ;
input E ;
input PRE ;
endmodule /* DFN0E1P0 */

module DFN0E1P1 (
  Q,
  CLK,
  D,
  E,
  PRE
)
;
output Q ;
input CLK ;
input D ;
input E ;
input PRE ;
endmodule /* DFN0E1P1 */

module DFN0P0 (
  Q,
  CLK,
  D,
  PRE
)
;
output Q ;
input CLK ;
input D ;
input PRE ;
endmodule /* DFN0P0 */

module DFN0P1 (
  Q,
  CLK,
  D,
  PRE
)
;
output Q ;
input CLK ;
input D ;
input PRE ;
endmodule /* DFN0P1 */

module DFN0P1C1 (
  Q,
  CLK,
  CLR,
  D,
  PRE
)
;
output Q ;
input CLK ;
input CLR ;
input D ;
input PRE ;
endmodule /* DFN0P1C1 */

module DFN1 (
  Q,
  CLK,
  D
)
;
output Q ;
input CLK ;
input D ;
endmodule /* DFN1 */

module DFN1C0 (
  Q,
  CLK,
  CLR,
  D
)
;
output Q ;
input CLK ;
input CLR ;
input D ;
endmodule /* DFN1C0 */

module DFN1C1 (
  Q,
  CLK,
  CLR,
  D
)
;
output Q ;
input CLK ;
input CLR ;
input D ;
endmodule /* DFN1C1 */

module DFN1E0 (
  Q,
  CLK,
  D,
  E
)
;
output Q ;
input CLK ;
input D ;
input E ;
endmodule /* DFN1E0 */

module DFN1E0C0 (
  Q,
  CLK,
  CLR,
  D,
  E
)
;
output Q ;
input CLK ;
input CLR ;
input D ;
input E ;
endmodule /* DFN1E0C0 */

module DFN1E0C1 (
  Q,
  CLK,
  CLR,
  D,
  E
)
;
output Q ;
input CLK ;
input CLR ;
input D ;
input E ;
endmodule /* DFN1E0C1 */

module DFN1E0P0 (
  Q,
  CLK,
  D,
  E,
  PRE
)
;
output Q ;
input CLK ;
input D ;
input E ;
input PRE ;
endmodule /* DFN1E0P0 */

module DFN1E0P1 (
  Q,
  CLK,
  D,
  E,
  PRE
)
;
output Q ;
input CLK ;
input D ;
input E ;
input PRE ;
endmodule /* DFN1E0P1 */

module DFN1E1 (
  Q,
  CLK,
  D,
  E
)
;
output Q ;
input CLK ;
input D ;
input E ;
endmodule /* DFN1E1 */

module DFN1E1C0 (
  Q,
  CLK,
  CLR,
  D,
  E
)
;
output Q ;
input CLK ;
input CLR ;
input D ;
input E ;
endmodule /* DFN1E1C0 */

module DFN1E1C1 (
  Q,
  CLK,
  CLR,
  D,
  E
)
;
output Q ;
input CLK ;
input CLR ;
input D ;
input E ;
endmodule /* DFN1E1C1 */

module DFN1E1P0 (
  Q,
  CLK,
  D,
  E,
  PRE
)
;
output Q ;
input CLK ;
input D ;
input E ;
input PRE ;
endmodule /* DFN1E1P0 */

module DFN1E1P1 (
  Q,
  CLK,
  D,
  E,
  PRE
)
;
output Q ;
input CLK ;
input D ;
input E ;
input PRE ;
endmodule /* DFN1E1P1 */

module DFN1P0 (
  Q,
  CLK,
  D,
  PRE
)
;
output Q ;
input CLK ;
input D ;
input PRE ;
endmodule /* DFN1P0 */

module DFN1P1 (
  Q,
  CLK,
  D,
  PRE
)
;
output Q ;
input CLK ;
input D ;
input PRE ;
endmodule /* DFN1P1 */

module DFN1P1C1 (
  Q,
  CLK,
  CLR,
  D,
  PRE
)
;
output Q ;
input CLK ;
input CLR ;
input D ;
input PRE ;
endmodule /* DFN1P1C1 */

module DLI0 (
  QN,
  D,
  G
)
;
output QN ;
input D ;
input G ;
endmodule /* DLI0 */

module DLI0C0 (
  QN,
  CLR,
  D,
  G
)
;
output QN ;
input CLR ;
input D ;
input G ;
endmodule /* DLI0C0 */

module DLI0C1 (
  QN,
  CLR,
  D,
  G
)
;
output QN ;
input CLR ;
input D ;
input G ;
endmodule /* DLI0C1 */

module DLI0P0 (
  QN,
  D,
  G,
  PRE
)
;
output QN ;
input D ;
input G ;
input PRE ;
endmodule /* DLI0P0 */

module DLI0P1 (
  QN,
  D,
  G,
  PRE
)
;
output QN ;
input D ;
input G ;
input PRE ;
endmodule /* DLI0P1 */

module DLI0P1C1 (
  QN,
  CLR,
  D,
  G,
  PRE
)
;
output QN ;
input CLR ;
input D ;
input G ;
input PRE ;
endmodule /* DLI0P1C1 */

module DLI1 (
  QN,
  D,
  G
)
;
output QN ;
input D ;
input G ;
endmodule /* DLI1 */

module DLI1C0 (
  QN,
  CLR,
  D,
  G
)
;
output QN ;
input CLR ;
input D ;
input G ;
endmodule /* DLI1C0 */

module DLI1C1 (
  QN,
  CLR,
  D,
  G
)
;
output QN ;
input CLR ;
input D ;
input G ;
endmodule /* DLI1C1 */

module DLI1P0 (
  QN,
  D,
  G,
  PRE
)
;
output QN ;
input D ;
input G ;
input PRE ;
endmodule /* DLI1P0 */

module DLI1P1 (
  QN,
  D,
  G,
  PRE
)
;
output QN ;
input D ;
input G ;
input PRE ;
endmodule /* DLI1P1 */

module DLI1P1C1 (
  QN,
  CLR,
  D,
  G,
  PRE
)
;
output QN ;
input CLR ;
input D ;
input G ;
input PRE ;
endmodule /* DLI1P1C1 */

module DLN0 (
  Q,
  D,
  G
)
;
output Q ;
input D ;
input G ;
endmodule /* DLN0 */

module DLN0C0 (
  Q,
  CLR,
  D,
  G
)
;
output Q ;
input CLR ;
input D ;
input G ;
endmodule /* DLN0C0 */

module DLN0C1 (
  Q,
  CLR,
  D,
  G
)
;
output Q ;
input CLR ;
input D ;
input G ;
endmodule /* DLN0C1 */

module DLN0P0 (
  Q,
  D,
  G,
  PRE
)
;
output Q ;
input D ;
input G ;
input PRE ;
endmodule /* DLN0P0 */

module DLN0P1 (
  Q,
  D,
  G,
  PRE
)
;
output Q ;
input D ;
input G ;
input PRE ;
endmodule /* DLN0P1 */

module DLN0P1C1 (
  Q,
  CLR,
  D,
  G,
  PRE
)
;
output Q ;
input CLR ;
input D ;
input G ;
input PRE ;
endmodule /* DLN0P1C1 */

module DLN1 (
  Q,
  D,
  G
)
;
output Q ;
input D ;
input G ;
endmodule /* DLN1 */

module DLN1C0 (
  Q,
  CLR,
  D,
  G
)
;
output Q ;
input CLR ;
input D ;
input G ;
endmodule /* DLN1C0 */

module DLN1C1 (
  Q,
  CLR,
  D,
  G
)
;
output Q ;
input CLR ;
input D ;
input G ;
endmodule /* DLN1C1 */

module DLN1P0 (
  Q,
  D,
  G,
  PRE
)
;
output Q ;
input D ;
input G ;
input PRE ;
endmodule /* DLN1P0 */

module DLN1P1 (
  Q,
  D,
  G,
  PRE
)
;
output Q ;
input D ;
input G ;
input PRE ;
endmodule /* DLN1P1 */

module DLN1P1C1 (
  Q,
  CLR,
  D,
  G,
  PRE
)
;
output Q ;
input CLR ;
input D ;
input G ;
input PRE ;
endmodule /* DLN1P1C1 */

module GND (
  Y
)
;
output Y ;
endmodule /* GND */

module INBUF_A (
  Y,
  PAD
)
;
output Y ;
input PAD ;
endmodule /* INBUF_A */

module INBUF_DA (
  Y,
  PAD
)
;
output Y ;
input PAD ;
endmodule /* INBUF_DA */

module INBUF (
  Y,
  PAD
)
;
output Y ;
input PAD ;
endmodule /* INBUF */

module INBUF_GTL25 (
  Y,
  PAD
)
;
output Y ;
input PAD ;
endmodule /* INBUF_GTL25 */

module INBUF_GTL33 (
  Y,
  PAD
)
;
output Y ;
input PAD ;
endmodule /* INBUF_GTL33 */

module INBUF_GTLP25 (
  Y,
  PAD
)
;
output Y ;
input PAD ;
endmodule /* INBUF_GTLP25 */

module INBUF_GTLP33 (
  Y,
  PAD
)
;
output Y ;
input PAD ;
endmodule /* INBUF_GTLP33 */

module INBUF_HSTL_I (
  Y,
  PAD
)
;
output Y ;
input PAD ;
endmodule /* INBUF_HSTL_I */

module INBUF_HSTL_II (
  Y,
  PAD
)
;
output Y ;
input PAD ;
endmodule /* INBUF_HSTL_II */

module INBUF_LVCMOS15 (
  Y,
  PAD
)
;
output Y ;
input PAD ;
endmodule /* INBUF_LVCMOS15 */

module INBUF_LVCMOS15D (
  Y,
  PAD
)
;
output Y ;
input PAD ;
endmodule /* INBUF_LVCMOS15D */

module INBUF_LVCMOS15U (
  Y,
  PAD
)
;
output Y ;
input PAD ;
endmodule /* INBUF_LVCMOS15U */

module INBUF_LVCMOS18 (
  Y,
  PAD
)
;
output Y ;
input PAD ;
endmodule /* INBUF_LVCMOS18 */

module INBUF_LVCMOS18D (
  Y,
  PAD
)
;
output Y ;
input PAD ;
endmodule /* INBUF_LVCMOS18D */

module INBUF_LVCMOS18U (
  Y,
  PAD
)
;
output Y ;
input PAD ;
endmodule /* INBUF_LVCMOS18U */

module INBUF_LVCMOS25 (
  Y,
  PAD
)
;
output Y ;
input PAD ;
endmodule /* INBUF_LVCMOS25 */

module INBUF_LVCMOS25D (
  Y,
  PAD
)
;
output Y ;
input PAD ;
endmodule /* INBUF_LVCMOS25D */

module INBUF_LVCMOS25U (
  Y,
  PAD
)
;
output Y ;
input PAD ;
endmodule /* INBUF_LVCMOS25U */

module INBUF_LVCMOS33 (
  Y,
  PAD
)
;
output Y ;
input PAD ;
endmodule /* INBUF_LVCMOS33 */

module INBUF_LVCMOS33D (
  Y,
  PAD
)
;
output Y ;
input PAD ;
endmodule /* INBUF_LVCMOS33D */

module INBUF_LVCMOS33U (
  Y,
  PAD
)
;
output Y ;
input PAD ;
endmodule /* INBUF_LVCMOS33U */

module INBUF_LVCMOS5 (
  Y,
  PAD
)
;
output Y ;
input PAD ;
endmodule /* INBUF_LVCMOS5 */

module INBUF_LVCMOS5D (
  Y,
  PAD
)
;
output Y ;
input PAD ;
endmodule /* INBUF_LVCMOS5D */

module INBUF_LVCMOS5U (
  Y,
  PAD
)
;
output Y ;
input PAD ;
endmodule /* INBUF_LVCMOS5U */

module INBUF_PCI (
  Y,
  PAD
)
;
output Y ;
input PAD ;
endmodule /* INBUF_PCI */

module INBUF_PCIX (
  Y,
  PAD
)
;
output Y ;
input PAD ;
endmodule /* INBUF_PCIX */

module INBUF_SSTL2_I (
  Y,
  PAD
)
;
output Y ;
input PAD ;
endmodule /* INBUF_SSTL2_I */

module INBUF_SSTL2_II (
  Y,
  PAD
)
;
output Y ;
input PAD ;
endmodule /* INBUF_SSTL2_II */

module INBUF_SSTL3_I (
  Y,
  PAD
)
;
output Y ;
input PAD ;
endmodule /* INBUF_SSTL3_I */

module INBUF_SSTL3_II (
  Y,
  PAD
)
;
output Y ;
input PAD ;
endmodule /* INBUF_SSTL3_II */

module INV (
  Y,
  A
)
;
output Y ;
input A ;
endmodule /* INV */

module INVD (
  Y,
  A
)
;
output Y ;
input A ;
endmodule /* INVD */

module IOBI_IB_OB_EB (
  DOUT,
  EOUT,
  Y,
  D,
  E,
  YIN
)
;
output DOUT ;
output EOUT ;
output Y ;
input D ;
input E ;
input YIN ;
endmodule /* IOBI_IB_OB_EB */

module IOBI_IB_OB_ER (
  DOUT,
  EOUT,
  Y,
  D,
  E,
  OCLK,
  YIN
)
;
output DOUT ;
output EOUT ;
output Y ;
input D ;
input E ;
input OCLK ;
input YIN ;
endmodule /* IOBI_IB_OB_ER */

module IOBI_IB_OB_ERC (
  DOUT,
  EOUT,
  Y,
  CLR,
  D,
  E,
  OCLK,
  YIN
)
;
output DOUT ;
output EOUT ;
output Y ;
input CLR ;
input D ;
input E ;
input OCLK ;
input YIN ;
endmodule /* IOBI_IB_OB_ERC */

module IOBI_IB_OB_ERE (
  DOUT,
  EOUT,
  Y,
  D,
  E,
  OCE,
  OCLK,
  YIN
)
;
output DOUT ;
output EOUT ;
output Y ;
input D ;
input E ;
input OCE ;
input OCLK ;
input YIN ;
endmodule /* IOBI_IB_OB_ERE */

module IOBI_IB_OB_EREC (
  DOUT,
  EOUT,
  Y,
  CLR,
  D,
  E,
  OCE,
  OCLK,
  YIN
)
;
output DOUT ;
output EOUT ;
output Y ;
input CLR ;
input D ;
input E ;
input OCE ;
input OCLK ;
input YIN ;
endmodule /* IOBI_IB_OB_EREC */

module IOBI_IB_OB_EREP (
  DOUT,
  EOUT,
  Y,
  D,
  E,
  OCE,
  OCLK,
  PRE,
  YIN
)
;
output DOUT ;
output EOUT ;
output Y ;
input D ;
input E ;
input OCE ;
input OCLK ;
input PRE ;
input YIN ;
endmodule /* IOBI_IB_OB_EREP */

module IOBI_IB_OB_ERP (
  DOUT,
  EOUT,
  Y,
  D,
  E,
  OCLK,
  PRE,
  YIN
)
;
output DOUT ;
output EOUT ;
output Y ;
input D ;
input E ;
input OCLK ;
input PRE ;
input YIN ;
endmodule /* IOBI_IB_OB_ERP */

module IOBI_IB_OR_EB (
  DOUT,
  EOUT,
  Y,
  D,
  E,
  OCLK,
  YIN
)
;
output DOUT ;
output EOUT ;
output Y ;
input D ;
input E ;
input OCLK ;
input YIN ;
endmodule /* IOBI_IB_OR_EB */

module IOBI_IB_OR_ER (
  DOUT,
  EOUT,
  Y,
  D,
  E,
  OCLK,
  YIN
)
;
output DOUT ;
output EOUT ;
output Y ;
input D ;
input E ;
input OCLK ;
input YIN ;
endmodule /* IOBI_IB_OR_ER */

module IOBI_IB_ORC_EB (
  DOUT,
  EOUT,
  Y,
  CLR,
  D,
  E,
  OCLK,
  YIN
)
;
output DOUT ;
output EOUT ;
output Y ;
input CLR ;
input D ;
input E ;
input OCLK ;
input YIN ;
endmodule /* IOBI_IB_ORC_EB */

module IOBI_IB_ORC_ERC (
  DOUT,
  EOUT,
  Y,
  CLR,
  D,
  E,
  OCLK,
  YIN
)
;
output DOUT ;
output EOUT ;
output Y ;
input CLR ;
input D ;
input E ;
input OCLK ;
input YIN ;
endmodule /* IOBI_IB_ORC_ERC */

module IOBI_IB_ORE_EB (
  DOUT,
  EOUT,
  Y,
  D,
  E,
  OCE,
  OCLK,
  YIN
)
;
output DOUT ;
output EOUT ;
output Y ;
input D ;
input E ;
input OCE ;
input OCLK ;
input YIN ;
endmodule /* IOBI_IB_ORE_EB */

module IOBI_IB_ORE_ERE (
  DOUT,
  EOUT,
  Y,
  D,
  E,
  OCE,
  OCLK,
  YIN
)
;
output DOUT ;
output EOUT ;
output Y ;
input D ;
input E ;
input OCE ;
input OCLK ;
input YIN ;
endmodule /* IOBI_IB_ORE_ERE */

module IOBI_IB_OREC_EB (
  DOUT,
  EOUT,
  Y,
  CLR,
  D,
  E,
  OCE,
  OCLK,
  YIN
)
;
output DOUT ;
output EOUT ;
output Y ;
input CLR ;
input D ;
input E ;
input OCE ;
input OCLK ;
input YIN ;
endmodule /* IOBI_IB_OREC_EB */

module IOBI_IB_OREC_EREC (
  DOUT,
  EOUT,
  Y,
  CLR,
  D,
  E,
  OCE,
  OCLK,
  YIN
)
;
output DOUT ;
output EOUT ;
output Y ;
input CLR ;
input D ;
input E ;
input OCE ;
input OCLK ;
input YIN ;
endmodule /* IOBI_IB_OREC_EREC */

module IOBI_IB_OREP_EB (
  DOUT,
  EOUT,
  Y,
  D,
  E,
  OCE,
  OCLK,
  PRE,
  YIN
)
;
output DOUT ;
output EOUT ;
output Y ;
input D ;
input E ;
input OCE ;
input OCLK ;
input PRE ;
input YIN ;
endmodule /* IOBI_IB_OREP_EB */

module IOBI_IB_OREP_EREP (
  DOUT,
  EOUT,
  Y,
  D,
  E,
  OCE,
  OCLK,
  PRE,
  YIN
)
;
output DOUT ;
output EOUT ;
output Y ;
input D ;
input E ;
input OCE ;
input OCLK ;
input PRE ;
input YIN ;
endmodule /* IOBI_IB_OREP_EREP */

module IOBI_IB_ORP_EB (
  DOUT,
  EOUT,
  Y,
  D,
  E,
  OCLK,
  PRE,
  YIN
)
;
output DOUT ;
output EOUT ;
output Y ;
input D ;
input E ;
input OCLK ;
input PRE ;
input YIN ;
endmodule /* IOBI_IB_ORP_EB */

module IOBI_IB_ORP_ERP (
  DOUT,
  EOUT,
  Y,
  D,
  E,
  OCLK,
  PRE,
  YIN
)
;
output DOUT ;
output EOUT ;
output Y ;
input D ;
input E ;
input OCLK ;
input PRE ;
input YIN ;
endmodule /* IOBI_IB_ORP_ERP */

module IOBI_IR_OB_EB (
  DOUT,
  EOUT,
  Y,
  D,
  E,
  ICLK,
  YIN
)
;
output DOUT ;
output EOUT ;
output Y ;
input D ;
input E ;
input ICLK ;
input YIN ;
endmodule /* IOBI_IR_OB_EB */

module IOBI_IR_OB_ER (
  DOUT,
  EOUT,
  Y,
  D,
  E,
  ICLK,
  OCLK,
  YIN
)
;
output DOUT ;
output EOUT ;
output Y ;
input D ;
input E ;
input ICLK ;
input OCLK ;
input YIN ;
endmodule /* IOBI_IR_OB_ER */

module IOBI_IR_OB_ERE (
  DOUT,
  EOUT,
  Y,
  D,
  E,
  ICLK,
  OCE,
  OCLK,
  YIN
)
;
output DOUT ;
output EOUT ;
output Y ;
input D ;
input E ;
input ICLK ;
input OCE ;
input OCLK ;
input YIN ;
endmodule /* IOBI_IR_OB_ERE */

module IOBI_IR_OR_EB (
  DOUT,
  EOUT,
  Y,
  D,
  E,
  ICLK,
  OCLK,
  YIN
)
;
output DOUT ;
output EOUT ;
output Y ;
input D ;
input E ;
input ICLK ;
input OCLK ;
input YIN ;
endmodule /* IOBI_IR_OR_EB */

module IOBI_IR_OR_ER (
  DOUT,
  EOUT,
  Y,
  D,
  E,
  ICLK,
  OCLK,
  YIN
)
;
output DOUT ;
output EOUT ;
output Y ;
input D ;
input E ;
input ICLK ;
input OCLK ;
input YIN ;
endmodule /* IOBI_IR_OR_ER */

module IOBI_IR_ORE_EB (
  DOUT,
  EOUT,
  Y,
  D,
  E,
  ICLK,
  OCE,
  OCLK,
  YIN
)
;
output DOUT ;
output EOUT ;
output Y ;
input D ;
input E ;
input ICLK ;
input OCE ;
input OCLK ;
input YIN ;
endmodule /* IOBI_IR_ORE_EB */

module IOBI_IR_ORE_ERE (
  DOUT,
  EOUT,
  Y,
  D,
  E,
  ICLK,
  OCE,
  OCLK,
  YIN
)
;
output DOUT ;
output EOUT ;
output Y ;
input D ;
input E ;
input ICLK ;
input OCE ;
input OCLK ;
input YIN ;
endmodule /* IOBI_IR_ORE_ERE */

module IOBI_IRC_OB_EB (
  DOUT,
  EOUT,
  Y,
  CLR,
  D,
  E,
  ICLK,
  YIN
)
;
output DOUT ;
output EOUT ;
output Y ;
input CLR ;
input D ;
input E ;
input ICLK ;
input YIN ;
endmodule /* IOBI_IRC_OB_EB */

module IOBI_IRC_OB_ERC (
  DOUT,
  EOUT,
  Y,
  CLR,
  D,
  E,
  ICLK,
  OCLK,
  YIN
)
;
output DOUT ;
output EOUT ;
output Y ;
input CLR ;
input D ;
input E ;
input ICLK ;
input OCLK ;
input YIN ;
endmodule /* IOBI_IRC_OB_ERC */

module IOBI_IRC_OB_EREC (
  DOUT,
  EOUT,
  Y,
  CLR,
  D,
  E,
  ICLK,
  OCE,
  OCLK,
  YIN
)
;
output DOUT ;
output EOUT ;
output Y ;
input CLR ;
input D ;
input E ;
input ICLK ;
input OCE ;
input OCLK ;
input YIN ;
endmodule /* IOBI_IRC_OB_EREC */

module IOBI_IRC_ORC_EB (
  DOUT,
  EOUT,
  Y,
  CLR,
  D,
  E,
  ICLK,
  OCLK,
  YIN
)
;
output DOUT ;
output EOUT ;
output Y ;
input CLR ;
input D ;
input E ;
input ICLK ;
input OCLK ;
input YIN ;
endmodule /* IOBI_IRC_ORC_EB */

module IOBI_IRC_ORC_ERC (
  DOUT,
  EOUT,
  Y,
  CLR,
  D,
  E,
  ICLK,
  OCLK,
  YIN
)
;
output DOUT ;
output EOUT ;
output Y ;
input CLR ;
input D ;
input E ;
input ICLK ;
input OCLK ;
input YIN ;
endmodule /* IOBI_IRC_ORC_ERC */

module IOBI_IRC_OREC_EB (
  DOUT,
  EOUT,
  Y,
  CLR,
  D,
  E,
  ICLK,
  OCE,
  OCLK,
  YIN
)
;
output DOUT ;
output EOUT ;
output Y ;
input CLR ;
input D ;
input E ;
input ICLK ;
input OCE ;
input OCLK ;
input YIN ;
endmodule /* IOBI_IRC_OREC_EB */

module IOBI_IRC_OREC_EREC (
  DOUT,
  EOUT,
  Y,
  CLR,
  D,
  E,
  ICLK,
  OCE,
  OCLK,
  YIN
)
;
output DOUT ;
output EOUT ;
output Y ;
input CLR ;
input D ;
input E ;
input ICLK ;
input OCE ;
input OCLK ;
input YIN ;
endmodule /* IOBI_IRC_OREC_EREC */

module IOBI_IRE_OB_EB (
  DOUT,
  EOUT,
  Y,
  D,
  E,
  ICE,
  ICLK,
  YIN
)
;
output DOUT ;
output EOUT ;
output Y ;
input D ;
input E ;
input ICE ;
input ICLK ;
input YIN ;
endmodule /* IOBI_IRE_OB_EB */

module IOBI_IRE_OB_ER (
  DOUT,
  EOUT,
  Y,
  D,
  E,
  ICE,
  ICLK,
  OCLK,
  YIN
)
;
output DOUT ;
output EOUT ;
output Y ;
input D ;
input E ;
input ICE ;
input ICLK ;
input OCLK ;
input YIN ;
endmodule /* IOBI_IRE_OB_ER */

module IOBI_IRE_OB_ERE (
  DOUT,
  EOUT,
  Y,
  D,
  E,
  ICE,
  ICLK,
  OCE,
  OCLK,
  YIN
)
;
output DOUT ;
output EOUT ;
output Y ;
input D ;
input E ;
input ICE ;
input ICLK ;
input OCE ;
input OCLK ;
input YIN ;
endmodule /* IOBI_IRE_OB_ERE */

module IOBI_IRE_OR_EB (
  DOUT,
  EOUT,
  Y,
  D,
  E,
  ICE,
  ICLK,
  OCLK,
  YIN
)
;
output DOUT ;
output EOUT ;
output Y ;
input D ;
input E ;
input ICE ;
input ICLK ;
input OCLK ;
input YIN ;
endmodule /* IOBI_IRE_OR_EB */

module IOBI_IRE_OR_ER (
  DOUT,
  EOUT,
  Y,
  D,
  E,
  ICE,
  ICLK,
  OCLK,
  YIN
)
;
output DOUT ;
output EOUT ;
output Y ;
input D ;
input E ;
input ICE ;
input ICLK ;
input OCLK ;
input YIN ;
endmodule /* IOBI_IRE_OR_ER */

module IOBI_IRE_ORE_EB (
  DOUT,
  EOUT,
  Y,
  D,
  E,
  ICE,
  ICLK,
  OCE,
  OCLK,
  YIN
)
;
output DOUT ;
output EOUT ;
output Y ;
input D ;
input E ;
input ICE ;
input ICLK ;
input OCE ;
input OCLK ;
input YIN ;
endmodule /* IOBI_IRE_ORE_EB */

module IOBI_IRE_ORE_ERE (
  DOUT,
  EOUT,
  Y,
  D,
  E,
  ICE,
  ICLK,
  OCE,
  OCLK,
  YIN
)
;
output DOUT ;
output EOUT ;
output Y ;
input D ;
input E ;
input ICE ;
input ICLK ;
input OCE ;
input OCLK ;
input YIN ;
endmodule /* IOBI_IRE_ORE_ERE */

module IOBI_IREC_OB_EB (
  DOUT,
  EOUT,
  Y,
  CLR,
  D,
  E,
  ICE,
  ICLK,
  YIN
)
;
output DOUT ;
output EOUT ;
output Y ;
input CLR ;
input D ;
input E ;
input ICE ;
input ICLK ;
input YIN ;
endmodule /* IOBI_IREC_OB_EB */

module IOBI_IREC_OB_ERC (
  DOUT,
  EOUT,
  Y,
  CLR,
  D,
  E,
  ICE,
  ICLK,
  OCLK,
  YIN
)
;
output DOUT ;
output EOUT ;
output Y ;
input CLR ;
input D ;
input E ;
input ICE ;
input ICLK ;
input OCLK ;
input YIN ;
endmodule /* IOBI_IREC_OB_ERC */

module IOBI_IREC_OB_EREC (
  DOUT,
  EOUT,
  Y,
  CLR,
  D,
  E,
  ICE,
  ICLK,
  OCE,
  OCLK,
  YIN
)
;
output DOUT ;
output EOUT ;
output Y ;
input CLR ;
input D ;
input E ;
input ICE ;
input ICLK ;
input OCE ;
input OCLK ;
input YIN ;
endmodule /* IOBI_IREC_OB_EREC */

module IOBI_IREC_ORC_EB (
  DOUT,
  EOUT,
  Y,
  CLR,
  D,
  E,
  ICE,
  ICLK,
  OCLK,
  YIN
)
;
output DOUT ;
output EOUT ;
output Y ;
input CLR ;
input D ;
input E ;
input ICE ;
input ICLK ;
input OCLK ;
input YIN ;
endmodule /* IOBI_IREC_ORC_EB */

module IOBI_IREC_ORC_ERC (
  DOUT,
  EOUT,
  Y,
  CLR,
  D,
  E,
  ICE,
  ICLK,
  OCLK,
  YIN
)
;
output DOUT ;
output EOUT ;
output Y ;
input CLR ;
input D ;
input E ;
input ICE ;
input ICLK ;
input OCLK ;
input YIN ;
endmodule /* IOBI_IREC_ORC_ERC */

module IOBI_IREC_OREC_EB (
  DOUT,
  EOUT,
  Y,
  CLR,
  D,
  E,
  ICE,
  ICLK,
  OCE,
  OCLK,
  YIN
)
;
output DOUT ;
output EOUT ;
output Y ;
input CLR ;
input D ;
input E ;
input ICE ;
input ICLK ;
input OCE ;
input OCLK ;
input YIN ;
endmodule /* IOBI_IREC_OREC_EB */

module IOBI_IREC_OREC_EREC (
  DOUT,
  EOUT,
  Y,
  CLR,
  D,
  E,
  ICE,
  ICLK,
  OCE,
  OCLK,
  YIN
)
;
output DOUT ;
output EOUT ;
output Y ;
input CLR ;
input D ;
input E ;
input ICE ;
input ICLK ;
input OCE ;
input OCLK ;
input YIN ;
endmodule /* IOBI_IREC_OREC_EREC */

module IOBI_IREP_OB_EB (
  DOUT,
  EOUT,
  Y,
  D,
  E,
  ICE,
  ICLK,
  PRE,
  YIN
)
;
output DOUT ;
output EOUT ;
output Y ;
input D ;
input E ;
input ICE ;
input ICLK ;
input PRE ;
input YIN ;
endmodule /* IOBI_IREP_OB_EB */

module IOBI_IREP_OB_EREP (
  DOUT,
  EOUT,
  Y,
  D,
  E,
  ICE,
  ICLK,
  OCE,
  OCLK,
  PRE,
  YIN
)
;
output DOUT ;
output EOUT ;
output Y ;
input D ;
input E ;
input ICE ;
input ICLK ;
input OCE ;
input OCLK ;
input PRE ;
input YIN ;
endmodule /* IOBI_IREP_OB_EREP */

module IOBI_IREP_OB_ERP (
  DOUT,
  EOUT,
  Y,
  D,
  E,
  ICE,
  ICLK,
  OCLK,
  PRE,
  YIN
)
;
output DOUT ;
output EOUT ;
output Y ;
input D ;
input E ;
input ICE ;
input ICLK ;
input OCLK ;
input PRE ;
input YIN ;
endmodule /* IOBI_IREP_OB_ERP */

module IOBI_IREP_OREP_EB (
  DOUT,
  EOUT,
  Y,
  D,
  E,
  ICE,
  ICLK,
  OCE,
  OCLK,
  PRE,
  YIN
)
;
output DOUT ;
output EOUT ;
output Y ;
input D ;
input E ;
input ICE ;
input ICLK ;
input OCE ;
input OCLK ;
input PRE ;
input YIN ;
endmodule /* IOBI_IREP_OREP_EB */

module IOBI_IREP_OREP_EREP (
  DOUT,
  EOUT,
  Y,
  D,
  E,
  ICE,
  ICLK,
  OCE,
  OCLK,
  PRE,
  YIN
)
;
output DOUT ;
output EOUT ;
output Y ;
input D ;
input E ;
input ICE ;
input ICLK ;
input OCE ;
input OCLK ;
input PRE ;
input YIN ;
endmodule /* IOBI_IREP_OREP_EREP */

module IOBI_IREP_ORP_EB (
  DOUT,
  EOUT,
  Y,
  D,
  E,
  ICE,
  ICLK,
  OCLK,
  PRE,
  YIN
)
;
output DOUT ;
output EOUT ;
output Y ;
input D ;
input E ;
input ICE ;
input ICLK ;
input OCLK ;
input PRE ;
input YIN ;
endmodule /* IOBI_IREP_ORP_EB */

module IOBI_IREP_ORP_ERP (
  DOUT,
  EOUT,
  Y,
  D,
  E,
  ICE,
  ICLK,
  OCLK,
  PRE,
  YIN
)
;
output DOUT ;
output EOUT ;
output Y ;
input D ;
input E ;
input ICE ;
input ICLK ;
input OCLK ;
input PRE ;
input YIN ;
endmodule /* IOBI_IREP_ORP_ERP */

module IOBI_IRP_OB_EB (
  DOUT,
  EOUT,
  Y,
  D,
  E,
  ICLK,
  PRE,
  YIN
)
;
output DOUT ;
output EOUT ;
output Y ;
input D ;
input E ;
input ICLK ;
input PRE ;
input YIN ;
endmodule /* IOBI_IRP_OB_EB */

module IOBI_IRP_OB_EREP (
  DOUT,
  EOUT,
  Y,
  D,
  E,
  ICLK,
  OCE,
  OCLK,
  PRE,
  YIN
)
;
output DOUT ;
output EOUT ;
output Y ;
input D ;
input E ;
input ICLK ;
input OCE ;
input OCLK ;
input PRE ;
input YIN ;
endmodule /* IOBI_IRP_OB_EREP */

module IOBI_IRP_OB_ERP (
  DOUT,
  EOUT,
  Y,
  D,
  E,
  ICLK,
  OCLK,
  PRE,
  YIN
)
;
output DOUT ;
output EOUT ;
output Y ;
input D ;
input E ;
input ICLK ;
input OCLK ;
input PRE ;
input YIN ;
endmodule /* IOBI_IRP_OB_ERP */

module IOBI_IRP_OREP_EB (
  DOUT,
  EOUT,
  Y,
  D,
  E,
  ICLK,
  OCE,
  OCLK,
  PRE,
  YIN
)
;
output DOUT ;
output EOUT ;
output Y ;
input D ;
input E ;
input ICLK ;
input OCE ;
input OCLK ;
input PRE ;
input YIN ;
endmodule /* IOBI_IRP_OREP_EB */

module IOBI_IRP_OREP_EREP (
  DOUT,
  EOUT,
  Y,
  D,
  E,
  ICLK,
  OCE,
  OCLK,
  PRE,
  YIN
)
;
output DOUT ;
output EOUT ;
output Y ;
input D ;
input E ;
input ICLK ;
input OCE ;
input OCLK ;
input PRE ;
input YIN ;
endmodule /* IOBI_IRP_OREP_EREP */

module IOBI_IRP_ORP_EB (
  DOUT,
  EOUT,
  Y,
  D,
  E,
  ICLK,
  OCLK,
  PRE,
  YIN
)
;
output DOUT ;
output EOUT ;
output Y ;
input D ;
input E ;
input ICLK ;
input OCLK ;
input PRE ;
input YIN ;
endmodule /* IOBI_IRP_ORP_EB */

module IOBI_IRP_ORP_ERP (
  DOUT,
  EOUT,
  Y,
  D,
  E,
  ICLK,
  OCLK,
  PRE,
  YIN
)
;
output DOUT ;
output EOUT ;
output Y ;
input D ;
input E ;
input ICLK ;
input OCLK ;
input PRE ;
input YIN ;
endmodule /* IOBI_IRP_ORP_ERP */

module IOIN_IB (
  Y,
  YIN
)
;
output Y ;
input YIN ;
endmodule /* IOIN_IB */

module IOIN_IR (
  Y,
  ICLK,
  YIN
)
;
output Y ;
input ICLK ;
input YIN ;
endmodule /* IOIN_IR */

module IOIN_IRC (
  Y,
  CLR,
  ICLK,
  YIN
)
;
output Y ;
input CLR ;
input ICLK ;
input YIN ;
endmodule /* IOIN_IRC */

module IOIN_IRE (
  Y,
  ICE,
  ICLK,
  YIN
)
;
output Y ;
input ICE ;
input ICLK ;
input YIN ;
endmodule /* IOIN_IRE */

module IOIN_IREC (
  Y,
  CLR,
  ICE,
  ICLK,
  YIN
)
;
output Y ;
input CLR ;
input ICE ;
input ICLK ;
input YIN ;
endmodule /* IOIN_IREC */

module IOIN_IREP (
  Y,
  ICE,
  ICLK,
  PRE,
  YIN
)
;
output Y ;
input ICE ;
input ICLK ;
input PRE ;
input YIN ;
endmodule /* IOIN_IREP */

module IOIN_IRP (
  Y,
  ICLK,
  PRE,
  YIN
)
;
output Y ;
input ICLK ;
input PRE ;
input YIN ;
endmodule /* IOIN_IRP */

module IOPAD_BI (
  PAD,
  Y,
  D,
  E
)
;
inout PAD /* synthesis syn_tristate = 1 */ ;
output Y ;
input D ;
input E ;
endmodule /* IOPAD_BI */

module IOPAD_BI_D (
  PAD,
  Y,
  D,
  E
)
;
inout PAD /* synthesis syn_tristate = 1 */ ;
output Y ;
input D ;
input E ;
endmodule /* IOPAD_BI_D */

module IOPAD_BI_U (
  PAD,
  Y,
  D,
  E
)
;
inout PAD /* synthesis syn_tristate = 1 */ ;
output Y ;
input D ;
input E ;
endmodule /* IOPAD_BI_U */

module IOPAD_IN (
  Y,
  PAD
)
;
output Y ;
input PAD ;
endmodule /* IOPAD_IN */

module IOPAD_IN_D (
  Y,
  PAD
)
;
output Y ;
input PAD ;
endmodule /* IOPAD_IN_D */

module IOPAD_IN_U (
  Y,
  PAD
)
;
output Y ;
input PAD ;
endmodule /* IOPAD_IN_U */

module IOPAD_A_IN (
  Y,
  PAD
)
;
output Y ;
input PAD ;
endmodule /* IOPAD_A_IN */

module IOPAD_DA_IN (
  Y,
  PAD
)
;
output Y ;
input PAD ;
endmodule /* IOPAD_DA_IN */

module IOPAD_TRI (
  PAD,
  D,
  E
)
;
output PAD /* synthesis syn_tristate = 1 */ ;
input D ;
input E ;
endmodule /* IOPAD_TRI */

module IOPAD_TRI_D (
  PAD,
  D,
  E
)
;
output PAD /* synthesis syn_tristate = 1 */ ;
input D ;
input E ;
endmodule /* IOPAD_TRI_D */

module IOPAD_TRI_U (
  PAD,
  D,
  E
)
;
output PAD /* synthesis syn_tristate = 1 */ ;
input D ;
input E ;
endmodule /* IOPAD_TRI_U */

module IOPADN_IN (
  N2POUT,
  PAD
)
;
output N2POUT ;
input PAD ;
endmodule /* IOPADN_IN */

module IOPADN_OUT (
  PAD,
  DB
)
;
output PAD ;
input DB ;
endmodule /* IOPADN_OUT */

module IOPAD_A_OUT (
  PAD,
  D
)
;
output PAD ;
input D ;
endmodule /* IOPAD_A_OUT */

module IOPADN_TRI (
  PAD,
  DB,
  E
)
;
output PAD /* synthesis syn_tristate = 1 */ ;
input DB ;
input E ;
endmodule /* IOPADN_TRI */

module IOPADP_BI (
  PAD,
  Y,
  D,
  E,
  N2PIN
)
;
inout PAD /* synthesis syn_tristate = 1 */ ;
output Y ;
input D ;
input E ;
input N2PIN ;
endmodule /* IOPADP_BI */

module IOPADN_BI (
  PAD,
  N2POUT,
  DB,
  E
)
;
inout PAD /* synthesis syn_tristate = 1 */ ;
output N2POUT ;
input DB ;
input E ;
endmodule /* IOPADN_BI */

module IOPADP_TRI (
  PAD,
  D,
  E
)
;
output PAD /* synthesis syn_tristate = 1 */ ;
input D ;
input E ;
endmodule /* IOPADP_TRI */

module IOTRI_OB_EB (
  DOUT,
  EOUT,
  D,
  E
)
;
output DOUT ;
output EOUT ;
input D ;
input E ;
endmodule /* IOTRI_OB_EB */

module IOTRI_OB_ER (
  DOUT,
  EOUT,
  D,
  E,
  OCLK
)
;
output DOUT ;
output EOUT ;
input D ;
input E ;
input OCLK ;
endmodule /* IOTRI_OB_ER */

module IOTRI_OB_ERC (
  DOUT,
  EOUT,
  CLR,
  D,
  E,
  OCLK
)
;
output DOUT ;
output EOUT ;
input CLR ;
input D ;
input E ;
input OCLK ;
endmodule /* IOTRI_OB_ERC */

module IOTRI_OB_ERE (
  DOUT,
  EOUT,
  D,
  E,
  OCE,
  OCLK
)
;
output DOUT ;
output EOUT ;
input D ;
input E ;
input OCE ;
input OCLK ;
endmodule /* IOTRI_OB_ERE */

module IOTRI_OB_EREC (
  DOUT,
  EOUT,
  CLR,
  D,
  E,
  OCE,
  OCLK
)
;
output DOUT ;
output EOUT ;
input CLR ;
input D ;
input E ;
input OCE ;
input OCLK ;
endmodule /* IOTRI_OB_EREC */

module IOTRI_OB_EREP (
  DOUT,
  EOUT,
  D,
  E,
  OCE,
  OCLK,
  PRE
)
;
output DOUT ;
output EOUT ;
input D ;
input E ;
input OCE ;
input OCLK ;
input PRE ;
endmodule /* IOTRI_OB_EREP */

module IOTRI_OB_ERP (
  DOUT,
  EOUT,
  D,
  E,
  OCLK,
  PRE
)
;
output DOUT ;
output EOUT ;
input D ;
input E ;
input OCLK ;
input PRE ;
endmodule /* IOTRI_OB_ERP */

module IOTRI_OR_EB (
  DOUT,
  EOUT,
  D,
  E,
  OCLK
)
;
output DOUT ;
output EOUT ;
input D ;
input E ;
input OCLK ;
endmodule /* IOTRI_OR_EB */

module IOTRI_OR_ER (
  DOUT,
  EOUT,
  D,
  E,
  OCLK
)
;
output DOUT ;
output EOUT ;
input D ;
input E ;
input OCLK ;
endmodule /* IOTRI_OR_ER */

module IOTRI_ORC_EB (
  DOUT,
  EOUT,
  CLR,
  D,
  E,
  OCLK
)
;
output DOUT ;
output EOUT ;
input CLR ;
input D ;
input E ;
input OCLK ;
endmodule /* IOTRI_ORC_EB */

module IOTRI_ORC_ERC (
  DOUT,
  EOUT,
  CLR,
  D,
  E,
  OCLK
)
;
output DOUT ;
output EOUT ;
input CLR ;
input D ;
input E ;
input OCLK ;
endmodule /* IOTRI_ORC_ERC */

module IOTRI_ORE_EB (
  DOUT,
  EOUT,
  D,
  E,
  OCE,
  OCLK
)
;
output DOUT ;
output EOUT ;
input D ;
input E ;
input OCE ;
input OCLK ;
endmodule /* IOTRI_ORE_EB */

module IOTRI_ORE_ERE (
  DOUT,
  EOUT,
  D,
  E,
  OCE,
  OCLK
)
;
output DOUT ;
output EOUT ;
input D ;
input E ;
input OCE ;
input OCLK ;
endmodule /* IOTRI_ORE_ERE */

module IOTRI_OREC_EB (
  DOUT,
  EOUT,
  CLR,
  D,
  E,
  OCE,
  OCLK
)
;
output DOUT ;
output EOUT ;
input CLR ;
input D ;
input E ;
input OCE ;
input OCLK ;
endmodule /* IOTRI_OREC_EB */

module IOTRI_OREC_EREC (
  DOUT,
  EOUT,
  CLR,
  D,
  E,
  OCE,
  OCLK
)
;
output DOUT ;
output EOUT ;
input CLR ;
input D ;
input E ;
input OCE ;
input OCLK ;
endmodule /* IOTRI_OREC_EREC */

module IOTRI_OREP_EB (
  DOUT,
  EOUT,
  D,
  E,
  OCE,
  OCLK,
  PRE
)
;
output DOUT ;
output EOUT ;
input D ;
input E ;
input OCE ;
input OCLK ;
input PRE ;
endmodule /* IOTRI_OREP_EB */

module IOTRI_OREP_EREP (
  DOUT,
  EOUT,
  D,
  E,
  OCE,
  OCLK,
  PRE
)
;
output DOUT ;
output EOUT ;
input D ;
input E ;
input OCE ;
input OCLK ;
input PRE ;
endmodule /* IOTRI_OREP_EREP */

module IOTRI_ORP_EB (
  DOUT,
  EOUT,
  D,
  E,
  OCLK,
  PRE
)
;
output DOUT ;
output EOUT ;
input D ;
input E ;
input OCLK ;
input PRE ;
endmodule /* IOTRI_ORP_EB */

module IOTRI_ORP_ERP (
  DOUT,
  EOUT,
  D,
  E,
  OCLK,
  PRE
)
;
output DOUT ;
output EOUT ;
input D ;
input E ;
input OCLK ;
input PRE ;
endmodule /* IOTRI_ORP_ERP */

module MAJ3 (
  Y,
  A,
  B,
  C
)
;
output Y ;
input A ;
input B ;
input C ;
endmodule /* MAJ3 */

module MAJ3X (
  Y,
  A,
  B,
  C
)
;
output Y ;
input A ;
input B ;
input C ;
endmodule /* MAJ3X */

module MAJ3XI (
  Y,
  A,
  B,
  C
)
;
output Y ;
input A ;
input B ;
input C ;
endmodule /* MAJ3XI */

module MIN3 (
  Y,
  A,
  B,
  C
)
;
output Y ;
input A ;
input B ;
input C ;
endmodule /* MIN3 */

module MIN3X (
  Y,
  A,
  B,
  C
)
;
output Y ;
input A ;
input B ;
input C ;
endmodule /* MIN3X */

module MIN3XI (
  Y,
  A,
  B,
  C
)
;
output Y ;
input A ;
input B ;
input C ;
endmodule /* MIN3XI */

module MX2 (
  Y,
  A,
  B,
  S
)
;
output Y ;
input A ;
input B ;
input S ;
endmodule /* MX2 */

module MX2A (
  Y,
  A,
  B,
  S
)
;
output Y ;
input A ;
input B ;
input S ;
endmodule /* MX2A */

module MX2B (
  Y,
  A,
  B,
  S
)
;
output Y ;
input A ;
input B ;
input S ;
endmodule /* MX2B */

module MX2C (
  Y,
  A,
  B,
  S
)
;
output Y ;
input A ;
input B ;
input S ;
endmodule /* MX2C */

module NAND2 (
  Y,
  A,
  B
)
;
output Y ;
input A ;
input B ;
endmodule /* NAND2 */

module NAND2A (
  Y,
  A,
  B
)
;
output Y ;
input A ;
input B ;
endmodule /* NAND2A */

module NAND2B (
  Y,
  A,
  B
)
;
output Y ;
input A ;
input B ;
endmodule /* NAND2B */

module NAND3 (
  Y,
  A,
  B,
  C
)
;
output Y ;
input A ;
input B ;
input C ;
endmodule /* NAND3 */

module NAND3A (
  Y,
  A,
  B,
  C
)
;
output Y ;
input A ;
input B ;
input C ;
endmodule /* NAND3A */

module NAND3B (
  Y,
  A,
  B,
  C
)
;
output Y ;
input A ;
input B ;
input C ;
endmodule /* NAND3B */

module NAND3C (
  Y,
  A,
  B,
  C
)
;
output Y ;
input A ;
input B ;
input C ;
endmodule /* NAND3C */

module NOR2 (
  Y,
  A,
  B
)
;
output Y ;
input A ;
input B ;
endmodule /* NOR2 */

module NOR2A (
  Y,
  A,
  B
)
;
output Y ;
input A ;
input B ;
endmodule /* NOR2A */

module NOR2B (
  Y,
  A,
  B
)
;
output Y ;
input A ;
input B ;
endmodule /* NOR2B */

module NOR3 (
  Y,
  A,
  B,
  C
)
;
output Y ;
input A ;
input B ;
input C ;
endmodule /* NOR3 */

module NOR3A (
  Y,
  A,
  B,
  C
)
;
output Y ;
input A ;
input B ;
input C ;
endmodule /* NOR3A */

module NOR3B (
  Y,
  A,
  B,
  C
)
;
output Y ;
input A ;
input B ;
input C ;
endmodule /* NOR3B */

module NOR3C (
  Y,
  A,
  B,
  C
)
;
output Y ;
input A ;
input B ;
input C ;
endmodule /* NOR3C */

module OA1 (
  Y,
  A,
  B,
  C
)
;
output Y ;
input A ;
input B ;
input C ;
endmodule /* OA1 */

module OA1A (
  Y,
  A,
  B,
  C
)
;
output Y ;
input A ;
input B ;
input C ;
endmodule /* OA1A */

module OA1B (
  Y,
  A,
  B,
  C
)
;
output Y ;
input A ;
input B ;
input C ;
endmodule /* OA1B */

module OA1C (
  Y,
  A,
  B,
  C
)
;
output Y ;
input A ;
input B ;
input C ;
endmodule /* OA1C */

module OAI1 (
  Y,
  A,
  B,
  C
)
;
output Y ;
input A ;
input B ;
input C ;
endmodule /* OAI1 */

module OR2 (
  Y,
  A,
  B
)
;
output Y ;
input A ;
input B ;
endmodule /* OR2 */

module OR2A (
  Y,
  A,
  B
)
;
output Y ;
input A ;
input B ;
endmodule /* OR2A */

module OR2B (
  Y,
  A,
  B
)
;
output Y ;
input A ;
input B ;
endmodule /* OR2B */

module OR3 (
  Y,
  A,
  B,
  C
)
;
output Y ;
input A ;
input B ;
input C ;
endmodule /* OR3 */

module OR3A (
  Y,
  A,
  B,
  C
)
;
output Y ;
input A ;
input B ;
input C ;
endmodule /* OR3A */

module OR3B (
  Y,
  A,
  B,
  C
)
;
output Y ;
input A ;
input B ;
input C ;
endmodule /* OR3B */

module OR3C (
  Y,
  A,
  B,
  C
)
;
output Y ;
input A ;
input B ;
input C ;
endmodule /* OR3C */

module OUTBUF_A (
  PAD,
  D
)
;
output PAD ;
input D ;
endmodule /* OUTBUF_A */

module OUTBUF (
  PAD,
  D
)
;
output PAD ;
input D ;
endmodule /* OUTBUF */

module OUTBUF_F_2 (
  PAD,
  D
)
;
output PAD ;
input D ;
endmodule /* OUTBUF_F_2 */

module OUTBUF_F_4 (
  PAD,
  D
)
;
output PAD ;
input D ;
endmodule /* OUTBUF_F_4 */

module OUTBUF_F_6 (
  PAD,
  D
)
;
output PAD ;
input D ;
endmodule /* OUTBUF_F_6 */

module OUTBUF_F_8 (
  PAD,
  D
)
;
output PAD ;
input D ;
endmodule /* OUTBUF_F_8 */

module OUTBUF_F_12 (
  PAD,
  D
)
;
output PAD ;
input D ;
endmodule /* OUTBUF_F_12 */

module OUTBUF_F_16 (
  PAD,
  D
)
;
output PAD ;
input D ;
endmodule /* OUTBUF_F_16 */

module OUTBUF_F_24 (
  PAD,
  D
)
;
output PAD ;
input D ;
endmodule /* OUTBUF_F_24 */

module OUTBUF_GTL25 (
  PAD,
  D
)
;
output PAD ;
input D ;
endmodule /* OUTBUF_GTL25 */

module OUTBUF_GTL33 (
  PAD,
  D
)
;
output PAD ;
input D ;
endmodule /* OUTBUF_GTL33 */

module OUTBUF_GTLP25 (
  PAD,
  D
)
;
output PAD ;
input D ;
endmodule /* OUTBUF_GTLP25 */

module OUTBUF_GTLP33 (
  PAD,
  D
)
;
output PAD ;
input D ;
endmodule /* OUTBUF_GTLP33 */

module OUTBUF_HSTL_I (
  PAD,
  D
)
;
output PAD ;
input D ;
endmodule /* OUTBUF_HSTL_I */

module OUTBUF_HSTL_II (
  PAD,
  D
)
;
output PAD ;
input D ;
endmodule /* OUTBUF_HSTL_II */

module OUTBUF_LVCMOS15 (
  PAD,
  D
)
;
output PAD ;
input D ;
endmodule /* OUTBUF_LVCMOS15 */

module OUTBUF_LVCMOS18 (
  PAD,
  D
)
;
output PAD ;
input D ;
endmodule /* OUTBUF_LVCMOS18 */

module OUTBUF_LVCMOS25 (
  PAD,
  D
)
;
output PAD ;
input D ;
endmodule /* OUTBUF_LVCMOS25 */

module OUTBUF_LVCMOS33 (
  PAD,
  D
)
;
output PAD ;
input D ;
endmodule /* OUTBUF_LVCMOS33 */

module OUTBUF_LVCMOS5 (
  PAD,
  D
)
;
output PAD ;
input D ;
endmodule /* OUTBUF_LVCMOS5 */

module OUTBUF_PCI (
  PAD,
  D
)
;
output PAD ;
input D ;
endmodule /* OUTBUF_PCI */

module OUTBUF_PCIX (
  PAD,
  D
)
;
output PAD ;
input D ;
endmodule /* OUTBUF_PCIX */

module OUTBUF_S_2 (
  PAD,
  D
)
;
output PAD ;
input D ;
endmodule /* OUTBUF_S_2 */

module OUTBUF_S_4 (
  PAD,
  D
)
;
output PAD ;
input D ;
endmodule /* OUTBUF_S_4 */

module OUTBUF_S_6 (
  PAD,
  D
)
;
output PAD ;
input D ;
endmodule /* OUTBUF_S_6 */

module OUTBUF_S_8 (
  PAD,
  D
)
;
output PAD ;
input D ;
endmodule /* OUTBUF_S_8 */

module OUTBUF_S_12 (
  PAD,
  D
)
;
output PAD ;
input D ;
endmodule /* OUTBUF_S_12 */

module OUTBUF_S_16 (
  PAD,
  D
)
;
output PAD ;
input D ;
endmodule /* OUTBUF_S_16 */

module OUTBUF_S_24 (
  PAD,
  D
)
;
output PAD ;
input D ;
endmodule /* OUTBUF_S_24 */

module OUTBUF_SSTL2_I (
  PAD,
  D
)
;
output PAD ;
input D ;
endmodule /* OUTBUF_SSTL2_I */

module OUTBUF_SSTL2_II (
  PAD,
  D
)
;
output PAD ;
input D ;
endmodule /* OUTBUF_SSTL2_II */

module OUTBUF_SSTL3_I (
  PAD,
  D
)
;
output PAD ;
input D ;
endmodule /* OUTBUF_SSTL3_I */

module OUTBUF_SSTL3_II (
  PAD,
  D
)
;
output PAD ;
input D ;
endmodule /* OUTBUF_SSTL3_II */

module TRIBUFF (
  PAD,
  D,
  E
)
;
output PAD /* synthesis syn_tristate = 1 */ ;
input D ;
input E ;
endmodule /* TRIBUFF */

module TRIBUFF_F_2 (
  PAD,
  D,
  E
)
;
output PAD /* synthesis syn_tristate = 1 */ ;
input D ;
input E ;
endmodule /* TRIBUFF_F_2 */

module TRIBUFF_F_2D (
  PAD,
  D,
  E
)
;
output PAD /* synthesis syn_tristate = 1 */ ;
input D ;
input E ;
endmodule /* TRIBUFF_F_2D */

module TRIBUFF_F_2U (
  PAD,
  D,
  E
)
;
output PAD /* synthesis syn_tristate = 1 */ ;
input D ;
input E ;
endmodule /* TRIBUFF_F_2U */

module TRIBUFF_F_4 (
  PAD,
  D,
  E
)
;
output PAD /* synthesis syn_tristate = 1 */ ;
input D ;
input E ;
endmodule /* TRIBUFF_F_4 */

module TRIBUFF_F_4D (
  PAD,
  D,
  E
)
;
output PAD /* synthesis syn_tristate = 1 */ ;
input D ;
input E ;
endmodule /* TRIBUFF_F_4D */

module TRIBUFF_F_4U (
  PAD,
  D,
  E
)
;
output PAD /* synthesis syn_tristate = 1 */ ;
input D ;
input E ;
endmodule /* TRIBUFF_F_4U */

module TRIBUFF_F_6 (
  PAD,
  D,
  E
)
;
output PAD /* synthesis syn_tristate = 1 */ ;
input D ;
input E ;
endmodule /* TRIBUFF_F_6 */

module TRIBUFF_F_6D (
  PAD,
  D,
  E
)
;
output PAD /* synthesis syn_tristate = 1 */ ;
input D ;
input E ;
endmodule /* TRIBUFF_F_6D */

module TRIBUFF_F_6U (
  PAD,
  D,
  E
)
;
output PAD /* synthesis syn_tristate = 1 */ ;
input D ;
input E ;
endmodule /* TRIBUFF_F_6U */

module TRIBUFF_F_8 (
  PAD,
  D,
  E
)
;
output PAD /* synthesis syn_tristate = 1 */ ;
input D ;
input E ;
endmodule /* TRIBUFF_F_8 */

module TRIBUFF_F_8D (
  PAD,
  D,
  E
)
;
output PAD /* synthesis syn_tristate = 1 */ ;
input D ;
input E ;
endmodule /* TRIBUFF_F_8D */

module TRIBUFF_F_8U (
  PAD,
  D,
  E
)
;
output PAD /* synthesis syn_tristate = 1 */ ;
input D ;
input E ;
endmodule /* TRIBUFF_F_8U */

module TRIBUFF_F_12 (
  PAD,
  D,
  E
)
;
output PAD /* synthesis syn_tristate = 1 */ ;
input D ;
input E ;
endmodule /* TRIBUFF_F_12 */

module TRIBUFF_F_12D (
  PAD,
  D,
  E
)
;
output PAD /* synthesis syn_tristate = 1 */ ;
input D ;
input E ;
endmodule /* TRIBUFF_F_12D */

module TRIBUFF_F_12U (
  PAD,
  D,
  E
)
;
output PAD /* synthesis syn_tristate = 1 */ ;
input D ;
input E ;
endmodule /* TRIBUFF_F_12U */

module TRIBUFF_F_16 (
  PAD,
  D,
  E
)
;
output PAD /* synthesis syn_tristate = 1 */ ;
input D ;
input E ;
endmodule /* TRIBUFF_F_16 */

module TRIBUFF_F_16D (
  PAD,
  D,
  E
)
;
output PAD /* synthesis syn_tristate = 1 */ ;
input D ;
input E ;
endmodule /* TRIBUFF_F_16D */

module TRIBUFF_F_16U (
  PAD,
  D,
  E
)
;
output PAD /* synthesis syn_tristate = 1 */ ;
input D ;
input E ;
endmodule /* TRIBUFF_F_16U */

module TRIBUFF_F_24 (
  PAD,
  D,
  E
)
;
output PAD /* synthesis syn_tristate = 1 */ ;
input D ;
input E ;
endmodule /* TRIBUFF_F_24 */

module TRIBUFF_F_24D (
  PAD,
  D,
  E
)
;
output PAD /* synthesis syn_tristate = 1 */ ;
input D ;
input E ;
endmodule /* TRIBUFF_F_24D */

module TRIBUFF_F_24U (
  PAD,
  D,
  E
)
;
output PAD /* synthesis syn_tristate = 1 */ ;
input D ;
input E ;
endmodule /* TRIBUFF_F_24U */

module TRIBUFF_GTL25 (
  PAD,
  D,
  E
)
;
output PAD /* synthesis syn_tristate = 1 */ ;
input D ;
input E ;
endmodule /* TRIBUFF_GTL25 */

module TRIBUFF_GTL33 (
  PAD,
  D,
  E
)
;
output PAD /* synthesis syn_tristate = 1 */ ;
input D ;
input E ;
endmodule /* TRIBUFF_GTL33 */

module TRIBUFF_GTLP25 (
  PAD,
  D,
  E
)
;
output PAD /* synthesis syn_tristate = 1 */ ;
input D ;
input E ;
endmodule /* TRIBUFF_GTLP25 */

module TRIBUFF_GTLP33 (
  PAD,
  D,
  E
)
;
output PAD /* synthesis syn_tristate = 1 */ ;
input D ;
input E ;
endmodule /* TRIBUFF_GTLP33 */

module TRIBUFF_HSTL_I (
  PAD,
  D,
  E
)
;
output PAD /* synthesis syn_tristate = 1 */ ;
input D ;
input E ;
endmodule /* TRIBUFF_HSTL_I */

module TRIBUFF_HSTL_II (
  PAD,
  D,
  E
)
;
output PAD /* synthesis syn_tristate = 1 */ ;
input D ;
input E ;
endmodule /* TRIBUFF_HSTL_II */

module TRIBUFF_LVCMOS15 (
  PAD,
  D,
  E
)
;
output PAD /* synthesis syn_tristate = 1 */ ;
input D ;
input E ;
endmodule /* TRIBUFF_LVCMOS15 */

module TRIBUFF_LVCMOS15D (
  PAD,
  D,
  E
)
;
output PAD /* synthesis syn_tristate = 1 */ ;
input D ;
input E ;
endmodule /* TRIBUFF_LVCMOS15D */

module TRIBUFF_LVCMOS15U (
  PAD,
  D,
  E
)
;
output PAD /* synthesis syn_tristate = 1 */ ;
input D ;
input E ;
endmodule /* TRIBUFF_LVCMOS15U */

module TRIBUFF_LVCMOS18 (
  PAD,
  D,
  E
)
;
output PAD /* synthesis syn_tristate = 1 */ ;
input D ;
input E ;
endmodule /* TRIBUFF_LVCMOS18 */

module TRIBUFF_LVCMOS18D (
  PAD,
  D,
  E
)
;
output PAD /* synthesis syn_tristate = 1 */ ;
input D ;
input E ;
endmodule /* TRIBUFF_LVCMOS18D */

module TRIBUFF_LVCMOS18U (
  PAD,
  D,
  E
)
;
output PAD /* synthesis syn_tristate = 1 */ ;
input D ;
input E ;
endmodule /* TRIBUFF_LVCMOS18U */

module TRIBUFF_LVCMOS25 (
  PAD,
  D,
  E
)
;
output PAD /* synthesis syn_tristate = 1 */ ;
input D ;
input E ;
endmodule /* TRIBUFF_LVCMOS25 */

module TRIBUFF_LVCMOS25D (
  PAD,
  D,
  E
)
;
output PAD /* synthesis syn_tristate = 1 */ ;
input D ;
input E ;
endmodule /* TRIBUFF_LVCMOS25D */

module TRIBUFF_LVCMOS25U (
  PAD,
  D,
  E
)
;
output PAD /* synthesis syn_tristate = 1 */ ;
input D ;
input E ;
endmodule /* TRIBUFF_LVCMOS25U */

module TRIBUFF_LVCMOS33 (
  PAD,
  D,
  E
)
;
output PAD /* synthesis syn_tristate = 1 */ ;
input D ;
input E ;
endmodule /* TRIBUFF_LVCMOS33 */

module TRIBUFF_LVCMOS33D (
  PAD,
  D,
  E
)
;
output PAD /* synthesis syn_tristate = 1 */ ;
input D ;
input E ;
endmodule /* TRIBUFF_LVCMOS33D */

module TRIBUFF_LVCMOS33U (
  PAD,
  D,
  E
)
;
output PAD /* synthesis syn_tristate = 1 */ ;
input D ;
input E ;
endmodule /* TRIBUFF_LVCMOS33U */

module TRIBUFF_LVCMOS5 (
  PAD,
  D,
  E
)
;
output PAD /* synthesis syn_tristate = 1 */ ;
input D ;
input E ;
endmodule /* TRIBUFF_LVCMOS5 */

module TRIBUFF_LVCMOS5D (
  PAD,
  D,
  E
)
;
output PAD /* synthesis syn_tristate = 1 */ ;
input D ;
input E ;
endmodule /* TRIBUFF_LVCMOS5D */

module TRIBUFF_LVCMOS5U (
  PAD,
  D,
  E
)
;
output PAD /* synthesis syn_tristate = 1 */ ;
input D ;
input E ;
endmodule /* TRIBUFF_LVCMOS5U */

module TRIBUFF_PCI (
  PAD,
  D,
  E
)
;
output PAD /* synthesis syn_tristate = 1 */ ;
input D ;
input E ;
endmodule /* TRIBUFF_PCI */

module TRIBUFF_PCIX (
  PAD,
  D,
  E
)
;
output PAD /* synthesis syn_tristate = 1 */ ;
input D ;
input E ;
endmodule /* TRIBUFF_PCIX */

module TRIBUFF_S_2 (
  PAD,
  D,
  E
)
;
output PAD /* synthesis syn_tristate = 1 */ ;
input D ;
input E ;
endmodule /* TRIBUFF_S_2 */

module TRIBUFF_S_2D (
  PAD,
  D,
  E
)
;
output PAD /* synthesis syn_tristate = 1 */ ;
input D ;
input E ;
endmodule /* TRIBUFF_S_2D */

module TRIBUFF_S_2U (
  PAD,
  D,
  E
)
;
output PAD /* synthesis syn_tristate = 1 */ ;
input D ;
input E ;
endmodule /* TRIBUFF_S_2U */

module TRIBUFF_S_4 (
  PAD,
  D,
  E
)
;
output PAD /* synthesis syn_tristate = 1 */ ;
input D ;
input E ;
endmodule /* TRIBUFF_S_4 */

module TRIBUFF_S_4D (
  PAD,
  D,
  E
)
;
output PAD /* synthesis syn_tristate = 1 */ ;
input D ;
input E ;
endmodule /* TRIBUFF_S_4D */

module TRIBUFF_S_4U (
  PAD,
  D,
  E
)
;
output PAD /* synthesis syn_tristate = 1 */ ;
input D ;
input E ;
endmodule /* TRIBUFF_S_4U */

module TRIBUFF_S_6 (
  PAD,
  D,
  E
)
;
output PAD /* synthesis syn_tristate = 1 */ ;
input D ;
input E ;
endmodule /* TRIBUFF_S_6 */

module TRIBUFF_S_6D (
  PAD,
  D,
  E
)
;
output PAD /* synthesis syn_tristate = 1 */ ;
input D ;
input E ;
endmodule /* TRIBUFF_S_6D */

module TRIBUFF_S_6U (
  PAD,
  D,
  E
)
;
output PAD /* synthesis syn_tristate = 1 */ ;
input D ;
input E ;
endmodule /* TRIBUFF_S_6U */

module TRIBUFF_S_8 (
  PAD,
  D,
  E
)
;
output PAD /* synthesis syn_tristate = 1 */ ;
input D ;
input E ;
endmodule /* TRIBUFF_S_8 */

module TRIBUFF_S_8D (
  PAD,
  D,
  E
)
;
output PAD /* synthesis syn_tristate = 1 */ ;
input D ;
input E ;
endmodule /* TRIBUFF_S_8D */

module TRIBUFF_S_8U (
  PAD,
  D,
  E
)
;
output PAD /* synthesis syn_tristate = 1 */ ;
input D ;
input E ;
endmodule /* TRIBUFF_S_8U */

module TRIBUFF_S_12 (
  PAD,
  D,
  E
)
;
output PAD /* synthesis syn_tristate = 1 */ ;
input D ;
input E ;
endmodule /* TRIBUFF_S_12 */

module TRIBUFF_S_12D (
  PAD,
  D,
  E
)
;
output PAD /* synthesis syn_tristate = 1 */ ;
input D ;
input E ;
endmodule /* TRIBUFF_S_12D */

module TRIBUFF_S_12U (
  PAD,
  D,
  E
)
;
output PAD /* synthesis syn_tristate = 1 */ ;
input D ;
input E ;
endmodule /* TRIBUFF_S_12U */

module TRIBUFF_S_16 (
  PAD,
  D,
  E
)
;
output PAD /* synthesis syn_tristate = 1 */ ;
input D ;
input E ;
endmodule /* TRIBUFF_S_16 */

module TRIBUFF_S_16D (
  PAD,
  D,
  E
)
;
output PAD /* synthesis syn_tristate = 1 */ ;
input D ;
input E ;
endmodule /* TRIBUFF_S_16D */

module TRIBUFF_S_16U (
  PAD,
  D,
  E
)
;
output PAD /* synthesis syn_tristate = 1 */ ;
input D ;
input E ;
endmodule /* TRIBUFF_S_16U */

module TRIBUFF_S_24 (
  PAD,
  D,
  E
)
;
output PAD /* synthesis syn_tristate = 1 */ ;
input D ;
input E ;
endmodule /* TRIBUFF_S_24 */

module TRIBUFF_S_24D (
  PAD,
  D,
  E
)
;
output PAD /* synthesis syn_tristate = 1 */ ;
input D ;
input E ;
endmodule /* TRIBUFF_S_24D */

module TRIBUFF_S_24U (
  PAD,
  D,
  E
)
;
output PAD /* synthesis syn_tristate = 1 */ ;
input D ;
input E ;
endmodule /* TRIBUFF_S_24U */

module TRIBUFF_SSTL2_I (
  PAD,
  D,
  E
)
;
output PAD /* synthesis syn_tristate = 1 */ ;
input D ;
input E ;
endmodule /* TRIBUFF_SSTL2_I */

module TRIBUFF_SSTL2_II (
  PAD,
  D,
  E
)
;
output PAD /* synthesis syn_tristate = 1 */ ;
input D ;
input E ;
endmodule /* TRIBUFF_SSTL2_II */

module TRIBUFF_SSTL3_I (
  PAD,
  D,
  E
)
;
output PAD /* synthesis syn_tristate = 1 */ ;
input D ;
input E ;
endmodule /* TRIBUFF_SSTL3_I */

module TRIBUFF_SSTL3_II (
  PAD,
  D,
  E
)
;
output PAD /* synthesis syn_tristate = 1 */ ;
input D ;
input E ;
endmodule /* TRIBUFF_SSTL3_II */

module TRIBUFF_LVDS (
  PADN,
  PADP,
  D,
  E
)
;
output PADN /* synthesis syn_tristate = 1 */ ;
output PADP /* synthesis syn_tristate = 1 */ ;
input D ;
input E ;
endmodule /* TRIBUFF_LVDS */

module VCC (
  Y
)
;
output Y ;
endmodule /* VCC */

module XA1 (
  Y,
  A,
  B,
  C
)
;
output Y ;
input A ;
input B ;
input C ;
endmodule /* XA1 */

module XA1A (
  Y,
  A,
  B,
  C
)
;
output Y ;
input A ;
input B ;
input C ;
endmodule /* XA1A */

module XA1B (
  Y,
  A,
  B,
  C
)
;
output Y ;
input A ;
input B ;
input C ;
endmodule /* XA1B */

module XA1C (
  Y,
  A,
  B,
  C
)
;
output Y ;
input A ;
input B ;
input C ;
endmodule /* XA1C */

module XAI1 (
  Y,
  A,
  B,
  C
)
;
output Y ;
input A ;
input B ;
input C ;
endmodule /* XAI1 */

module XAI1A (
  Y,
  A,
  B,
  C
)
;
output Y ;
input A ;
input B ;
input C ;
endmodule /* XAI1A */

module XNOR2 (
  Y,
  A,
  B
)
;
output Y ;
input A ;
input B ;
endmodule /* XNOR2 */

module XNOR3 (
  Y,
  A,
  B,
  C
)
;
output Y ;
input A ;
input B ;
input C ;
endmodule /* XNOR3 */

module XO1 (
  Y,
  A,
  B,
  C
)
;
output Y ;
input A ;
input B ;
input C ;
endmodule /* XO1 */

module XO1A (
  Y,
  A,
  B,
  C
)
;
output Y ;
input A ;
input B ;
input C ;
endmodule /* XO1A */

module XOR2 (
  Y,
  A,
  B
)
;
output Y ;
input A ;
input B ;
endmodule /* XOR2 */

module XOR3 (
  Y,
  A,
  B,
  C
)
;
output Y ;
input A ;
input B ;
input C ;
endmodule /* XOR3 */

module ZOR3 (
  Y,
  A,
  B,
  C
)
;
output Y ;
input A ;
input B ;
input C ;
endmodule /* ZOR3 */

module ZOR3I (
  Y,
  A,
  B,
  C
)
;
output Y ;
input A ;
input B ;
input C ;
endmodule /* ZOR3I */

module CLKDLY (
  GL,
  CLK,
  DLYGL0,
  DLYGL1,
  DLYGL2,
  DLYGL3,
  DLYGL4
)
;
output GL ;
input CLK ;
input DLYGL0 ;
input DLYGL1 ;
input DLYGL2 ;
input DLYGL3 ;
input DLYGL4 ;
endmodule /* CLKDLY */

module CLKSRC (
  Y,
  A
)
;
output Y ;
input A ;
endmodule /* CLKSRC */

module CLKDIV_SDF (
  GL,
  CLK,
  ODIV0,
  ODIV1,
  ODIV2,
  ODIV3,
  ODIV4,
  ODIVHALF,
  RESET
)
;
output GL ;
input CLK ;
input ODIV0 ;
input ODIV1 ;
input ODIV2 ;
input ODIV3 ;
input ODIV4 ;
input ODIVHALF ;
input RESET ;
endmodule /* CLKDIV_SDF */

module CLKDLY_SDF (
  GL,
  CLK,
  DLYGL0,
  DLYGL1,
  DLYGL2,
  DLYGL3,
  DLYGL4
)
;
output GL ;
input CLK ;
input DLYGL0 ;
input DLYGL1 ;
input DLYGL2 ;
input DLYGL3 ;
input DLYGL4 ;
endmodule /* CLKDLY_SDF */

module CLKDIVDLY_SDF (
  GL,
  CLK,
  DLYGL0,
  DLYGL1,
  DLYGL2,
  DLYGL3,
  DLYGL4
)
;
output GL ;
input CLK ;
input DLYGL0 ;
input DLYGL1 ;
input DLYGL2 ;
input DLYGL3 ;
input DLYGL4 ;
endmodule /* CLKDIVDLY_SDF */

module CLKDIVDLY1_SDF (
  GL,
  Y,
  CLK,
  DLYGL0,
  DLYGL1,
  DLYGL2,
  DLYGL3,
  DLYGL4,
  DLYY0,
  DLYY1,
  DLYY2,
  DLYY3,
  DLYY4
)
;
output GL ;
output Y ;
input CLK ;
input DLYGL0 ;
input DLYGL1 ;
input DLYGL2 ;
input DLYGL3 ;
input DLYGL4 ;
input DLYY0 ;
input DLYY1 ;
input DLYY2 ;
input DLYY3 ;
input DLYY4 ;
endmodule /* CLKDIVDLY1_SDF */

module RCOSC (
  CLKOUT
)
;
output CLKOUT ;
endmodule /* RCOSC */

module DDR_OUT (
  Q,
  CLK,
  CLR,
  DF,
  DR
)
;
output Q ;
input CLK ;
input CLR ;
input DF ;
input DR ;
endmodule /* DDR_OUT */

module DDR_REG (
  QF,
  QR,
  CLK,
  CLR,
  D
)
;
output QF ;
output QR ;
input CLK ;
input CLR ;
input D ;
endmodule /* DDR_REG */

module FIFO4K18 (
  AEMPTY,
  AFULL,
  EMPTY,
  FULL,
  RD0,
  RD1,
  RD2,
  RD3,
  RD4,
  RD5,
  RD6,
  RD7,
  RD8,
  RD9,
  RD10,
  RD11,
  RD12,
  RD13,
  RD14,
  RD15,
  RD16,
  RD17,
  AEVAL11,
  AEVAL10,
  AEVAL9,
  AEVAL8,
  AEVAL7,
  AEVAL6,
  AEVAL5,
  AEVAL4,
  AEVAL3,
  AEVAL2,
  AEVAL1,
  AEVAL0,
  AFVAL11,
  AFVAL10,
  AFVAL9,
  AFVAL8,
  AFVAL7,
  AFVAL6,
  AFVAL5,
  AFVAL4,
  AFVAL3,
  AFVAL2,
  AFVAL1,
  AFVAL0,
  ESTOP,
  FSTOP,
  RCLK,
  REN,
  RBLK,
  RESET,
  RPIPE,
  RW2,
  RW1,
  RW0,
  WCLK,
  WD0,
  WD1,
  WD2,
  WD3,
  WD4,
  WD5,
  WD6,
  WD7,
  WD8,
  WD9,
  WD10,
  WD11,
  WD12,
  WD13,
  WD14,
  WD15,
  WD16,
  WD17,
  WEN,
  WBLK,
  WW2,
  WW1,
  WW0
)
;
output AEMPTY ;
output AFULL ;
output EMPTY ;
output FULL ;
output RD0 ;
output RD1 ;
output RD2 ;
output RD3 ;
output RD4 ;
output RD5 ;
output RD6 ;
output RD7 ;
output RD8 ;
output RD9 ;
output RD10 ;
output RD11 ;
output RD12 ;
output RD13 ;
output RD14 ;
output RD15 ;
output RD16 ;
output RD17 ;
input AEVAL11 ;
input AEVAL10 ;
input AEVAL9 ;
input AEVAL8 ;
input AEVAL7 ;
input AEVAL6 ;
input AEVAL5 ;
input AEVAL4 ;
input AEVAL3 ;
input AEVAL2 ;
input AEVAL1 ;
input AEVAL0 ;
input AFVAL11 ;
input AFVAL10 ;
input AFVAL9 ;
input AFVAL8 ;
input AFVAL7 ;
input AFVAL6 ;
input AFVAL5 ;
input AFVAL4 ;
input AFVAL3 ;
input AFVAL2 ;
input AFVAL1 ;
input AFVAL0 ;
input ESTOP ;
input FSTOP ;
input RCLK ;
input REN ;
input RBLK ;
input RESET ;
input RPIPE ;
input RW2 ;
input RW1 ;
input RW0 ;
input WCLK ;
input WD0 ;
input WD1 ;
input WD2 ;
input WD3 ;
input WD4 ;
input WD5 ;
input WD6 ;
input WD7 ;
input WD8 ;
input WD9 ;
input WD10 ;
input WD11 ;
input WD12 ;
input WD13 ;
input WD14 ;
input WD15 ;
input WD16 ;
input WD17 ;
input WEN ;
input WBLK ;
input WW2 ;
input WW1 ;
input WW0 ;
endmodule /* FIFO4K18 */

module PLLINT (
  Y,
  A
)
;
output Y ;
input A ;
endmodule /* PLLINT */

module RAM4K9 (
  DOUTA0,
  DOUTA1,
  DOUTA2,
  DOUTA3,
  DOUTA4,
  DOUTA5,
  DOUTA6,
  DOUTA7,
  DOUTA8,
  DOUTB0,
  DOUTB1,
  DOUTB2,
  DOUTB3,
  DOUTB4,
  DOUTB5,
  DOUTB6,
  DOUTB7,
  DOUTB8,
  ADDRA0,
  ADDRA1,
  ADDRA2,
  ADDRA3,
  ADDRA4,
  ADDRA5,
  ADDRA6,
  ADDRA7,
  ADDRA8,
  ADDRA9,
  ADDRA10,
  ADDRA11,
  ADDRB0,
  ADDRB1,
  ADDRB2,
  ADDRB3,
  ADDRB4,
  ADDRB5,
  ADDRB6,
  ADDRB7,
  ADDRB8,
  ADDRB9,
  ADDRB10,
  ADDRB11,
  BLKA,
  BLKB,
  CLKA,
  CLKB,
  DINA0,
  DINA1,
  DINA2,
  DINA3,
  DINA4,
  DINA5,
  DINA6,
  DINA7,
  DINA8,
  DINB0,
  DINB1,
  DINB2,
  DINB3,
  DINB4,
  DINB5,
  DINB6,
  DINB7,
  DINB8,
  PIPEA,
  PIPEB,
  RESET,
  WENA,
  WENB,
  WIDTHA1,
  WIDTHA0,
  WIDTHB1,
  WIDTHB0,
  WMODEA,
  WMODEB
)
;
output DOUTA0 ;
output DOUTA1 ;
output DOUTA2 ;
output DOUTA3 ;
output DOUTA4 ;
output DOUTA5 ;
output DOUTA6 ;
output DOUTA7 ;
output DOUTA8 ;
output DOUTB0 ;
output DOUTB1 ;
output DOUTB2 ;
output DOUTB3 ;
output DOUTB4 ;
output DOUTB5 ;
output DOUTB6 ;
output DOUTB7 ;
output DOUTB8 ;
input ADDRA0 ;
input ADDRA1 ;
input ADDRA2 ;
input ADDRA3 ;
input ADDRA4 ;
input ADDRA5 ;
input ADDRA6 ;
input ADDRA7 ;
input ADDRA8 ;
input ADDRA9 ;
input ADDRA10 ;
input ADDRA11 ;
input ADDRB0 ;
input ADDRB1 ;
input ADDRB2 ;
input ADDRB3 ;
input ADDRB4 ;
input ADDRB5 ;
input ADDRB6 ;
input ADDRB7 ;
input ADDRB8 ;
input ADDRB9 ;
input ADDRB10 ;
input ADDRB11 ;
input BLKA ;
input BLKB ;
input CLKA ;
input CLKB ;
input DINA0 ;
input DINA1 ;
input DINA2 ;
input DINA3 ;
input DINA4 ;
input DINA5 ;
input DINA6 ;
input DINA7 ;
input DINA8 ;
input DINB0 ;
input DINB1 ;
input DINB2 ;
input DINB3 ;
input DINB4 ;
input DINB5 ;
input DINB6 ;
input DINB7 ;
input DINB8 ;
input PIPEA ;
input PIPEB ;
input RESET ;
input WENA ;
input WENB ;
input WIDTHA1 ;
input WIDTHA0 ;
input WIDTHB1 ;
input WIDTHB0 ;
input WMODEA ;
input WMODEB ;
endmodule /* RAM4K9 */

module RAM512X18 (
  RD0,
  RD1,
  RD2,
  RD3,
  RD4,
  RD5,
  RD6,
  RD7,
  RD8,
  RD9,
  RD10,
  RD11,
  RD12,
  RD13,
  RD14,
  RD15,
  RD16,
  RD17,
  PIPE,
  RADDR0,
  RADDR1,
  RADDR2,
  RADDR3,
  RADDR4,
  RADDR5,
  RADDR6,
  RADDR7,
  RADDR8,
  RCLK,
  REN,
  RESET,
  RW1,
  RW0,
  WADDR0,
  WADDR1,
  WADDR2,
  WADDR3,
  WADDR4,
  WADDR5,
  WADDR6,
  WADDR7,
  WADDR8,
  WCLK,
  WD0,
  WD1,
  WD2,
  WD3,
  WD4,
  WD5,
  WD6,
  WD7,
  WD8,
  WD9,
  WD10,
  WD11,
  WD12,
  WD13,
  WD14,
  WD15,
  WD16,
  WD17,
  WEN,
  WW1,
  WW0
)
;
output RD0 ;
output RD1 ;
output RD2 ;
output RD3 ;
output RD4 ;
output RD5 ;
output RD6 ;
output RD7 ;
output RD8 ;
output RD9 ;
output RD10 ;
output RD11 ;
output RD12 ;
output RD13 ;
output RD14 ;
output RD15 ;
output RD16 ;
output RD17 ;
input PIPE ;
input RADDR0 ;
input RADDR1 ;
input RADDR2 ;
input RADDR3 ;
input RADDR4 ;
input RADDR5 ;
input RADDR6 ;
input RADDR7 ;
input RADDR8 ;
input RCLK ;
input REN ;
input RESET ;
input RW1 ;
input RW0 ;
input WADDR0 ;
input WADDR1 ;
input WADDR2 ;
input WADDR3 ;
input WADDR4 ;
input WADDR5 ;
input WADDR6 ;
input WADDR7 ;
input WADDR8 ;
input WCLK ;
input WD0 ;
input WD1 ;
input WD2 ;
input WD3 ;
input WD4 ;
input WD5 ;
input WD6 ;
input WD7 ;
input WD8 ;
input WD9 ;
input WD10 ;
input WD11 ;
input WD12 ;
input WD13 ;
input WD14 ;
input WD15 ;
input WD16 ;
input WD17 ;
input WEN ;
input WW1 ;
input WW0 ;
endmodule /* RAM512X18 */

module FLEXRAM4K9 (
  DOUTA0,
  DOUTA1,
  DOUTA2,
  DOUTA3,
  DOUTA4,
  DOUTA5,
  DOUTA6,
  DOUTA7,
  DOUTA8,
  DOUTB0,
  DOUTB1,
  DOUTB2,
  DOUTB3,
  DOUTB4,
  DOUTB5,
  DOUTB6,
  DOUTB7,
  DOUTB8,
  ADDRA0,
  ADDRA1,
  ADDRA2,
  ADDRA3,
  ADDRA4,
  ADDRA5,
  ADDRA6,
  ADDRA7,
  ADDRA8,
  ADDRA9,
  ADDRA10,
  ADDRA11,
  ADDRB0,
  ADDRB1,
  ADDRB2,
  ADDRB3,
  ADDRB4,
  ADDRB5,
  ADDRB6,
  ADDRB7,
  ADDRB8,
  ADDRB9,
  ADDRB10,
  ADDRB11,
  BLKA,
  BLKB,
  CLKA,
  CLKB,
  DINA0,
  DINA1,
  DINA2,
  DINA3,
  DINA4,
  DINA5,
  DINA6,
  DINA7,
  DINA8,
  DINB0,
  DINB1,
  DINB2,
  DINB3,
  DINB4,
  DINB5,
  DINB6,
  DINB7,
  DINB8,
  PIPEA,
  PIPEB,
  RESET,
  WENA,
  WENB,
  WIDTHA1,
  WIDTHA0,
  WIDTHB1,
  WIDTHB0,
  WMODEA,
  WMODEB
)
;
output DOUTA0 ;
output DOUTA1 ;
output DOUTA2 ;
output DOUTA3 ;
output DOUTA4 ;
output DOUTA5 ;
output DOUTA6 ;
output DOUTA7 ;
output DOUTA8 ;
output DOUTB0 ;
output DOUTB1 ;
output DOUTB2 ;
output DOUTB3 ;
output DOUTB4 ;
output DOUTB5 ;
output DOUTB6 ;
output DOUTB7 ;
output DOUTB8 ;
input ADDRA0 ;
input ADDRA1 ;
input ADDRA2 ;
input ADDRA3 ;
input ADDRA4 ;
input ADDRA5 ;
input ADDRA6 ;
input ADDRA7 ;
input ADDRA8 ;
input ADDRA9 ;
input ADDRA10 ;
input ADDRA11 ;
input ADDRB0 ;
input ADDRB1 ;
input ADDRB2 ;
input ADDRB3 ;
input ADDRB4 ;
input ADDRB5 ;
input ADDRB6 ;
input ADDRB7 ;
input ADDRB8 ;
input ADDRB9 ;
input ADDRB10 ;
input ADDRB11 ;
input BLKA ;
input BLKB ;
input CLKA ;
input CLKB ;
input DINA0 ;
input DINA1 ;
input DINA2 ;
input DINA3 ;
input DINA4 ;
input DINA5 ;
input DINA6 ;
input DINA7 ;
input DINA8 ;
input DINB0 ;
input DINB1 ;
input DINB2 ;
input DINB3 ;
input DINB4 ;
input DINB5 ;
input DINB6 ;
input DINB7 ;
input DINB8 ;
input PIPEA ;
input PIPEB ;
input RESET ;
input WENA ;
input WENB ;
input WIDTHA1 ;
input WIDTHA0 ;
input WIDTHB1 ;
input WIDTHB0 ;
input WMODEA ;
input WMODEB ;
endmodule /* FLEXRAM4K9 */

module FLEXRAM512X18 (
  RD0,
  RD1,
  RD2,
  RD3,
  RD4,
  RD5,
  RD6,
  RD7,
  RD8,
  RD9,
  RD10,
  RD11,
  RD12,
  RD13,
  RD14,
  RD15,
  RD16,
  RD17,
  PIPE,
  RADDR0,
  RADDR1,
  RADDR2,
  RADDR3,
  RADDR4,
  RADDR5,
  RADDR6,
  RADDR7,
  RADDR8,
  RCLK,
  REN,
  RESET,
  RW1,
  RW0,
  WADDR0,
  WADDR1,
  WADDR2,
  WADDR3,
  WADDR4,
  WADDR5,
  WADDR6,
  WADDR7,
  WADDR8,
  WCLK,
  WD0,
  WD1,
  WD2,
  WD3,
  WD4,
  WD5,
  WD6,
  WD7,
  WD8,
  WD9,
  WD10,
  WD11,
  WD12,
  WD13,
  WD14,
  WD15,
  WD16,
  WD17,
  WEN,
  WW1,
  WW0
)
;
output RD0 ;
output RD1 ;
output RD2 ;
output RD3 ;
output RD4 ;
output RD5 ;
output RD6 ;
output RD7 ;
output RD8 ;
output RD9 ;
output RD10 ;
output RD11 ;
output RD12 ;
output RD13 ;
output RD14 ;
output RD15 ;
output RD16 ;
output RD17 ;
input PIPE ;
input RADDR0 ;
input RADDR1 ;
input RADDR2 ;
input RADDR3 ;
input RADDR4 ;
input RADDR5 ;
input RADDR6 ;
input RADDR7 ;
input RADDR8 ;
input RCLK ;
input REN ;
input RESET ;
input RW1 ;
input RW0 ;
input WADDR0 ;
input WADDR1 ;
input WADDR2 ;
input WADDR3 ;
input WADDR4 ;
input WADDR5 ;
input WADDR6 ;
input WADDR7 ;
input WADDR8 ;
input WCLK ;
input WD0 ;
input WD1 ;
input WD2 ;
input WD3 ;
input WD4 ;
input WD5 ;
input WD6 ;
input WD7 ;
input WD8 ;
input WD9 ;
input WD10 ;
input WD11 ;
input WD12 ;
input WD13 ;
input WD14 ;
input WD15 ;
input WD16 ;
input WD17 ;
input WEN ;
input WW1 ;
input WW0 ;
endmodule /* FLEXRAM512X18 */

module UJTAG (
  TDO,
  UDRCAP,
  UDRCK,
  UDRSH,
  UDRUPD,
  UIREG0,
  UIREG1,
  UIREG2,
  UIREG3,
  UIREG4,
  UIREG5,
  UIREG6,
  UIREG7,
  URSTB,
  UTDI,
  TCK,
  TDI,
  TMS,
  TRSTB,
  UTDO
)
;
output TDO ;
output UDRCAP ;
output UDRCK ;
output UDRSH ;
output UDRUPD ;
output UIREG0 ;
output UIREG1 ;
output UIREG2 ;
output UIREG3 ;
output UIREG4 ;
output UIREG5 ;
output UIREG6 ;
output UIREG7 ;
output URSTB ;
output UTDI ;
input TCK ;
input TDI ;
input TMS ;
input TRSTB ;
input UTDO ;
endmodule /* UJTAG */

module IOBI_ID_OB_EB (
  DOUT,
  EOUT,
  YF,
  YR,
  CLR,
  D,
  E,
  ICLK,
  YIN
)
;
output DOUT ;
output EOUT ;
output YF ;
output YR ;
input CLR ;
input D ;
input E ;
input ICLK ;
input YIN ;
endmodule /* IOBI_ID_OB_EB */

module IOBI_IB_OD_EB (
  DOUT,
  EOUT,
  Y,
  CLR,
  DF,
  DR,
  E,
  OCLK,
  YIN
)
;
output DOUT ;
output EOUT ;
output Y ;
input CLR ;
input DF ;
input DR ;
input E ;
input OCLK ;
input YIN ;
endmodule /* IOBI_IB_OD_EB */

module IOBI_ID_OD_EB (
  DOUT,
  EOUT,
  YF,
  YR,
  CLR,
  DF,
  DR,
  E,
  ICLK,
  OCLK,
  YIN
)
;
output DOUT ;
output EOUT ;
output YF ;
output YR ;
input CLR ;
input DF ;
input DR ;
input E ;
input ICLK ;
input OCLK ;
input YIN ;
endmodule /* IOBI_ID_OD_EB */

module IOBI_ID_OD_ERC (
  DOUT,
  EOUT,
  YF,
  YR,
  CLR,
  DF,
  DR,
  E,
  ICLK,
  OCLK,
  YIN
)
;
output DOUT ;
output EOUT ;
output YF ;
output YR ;
input CLR ;
input DF ;
input DR ;
input E ;
input ICLK ;
input OCLK ;
input YIN ;
endmodule /* IOBI_ID_OD_ERC */

module IOIN_ID (
  YF,
  YR,
  CLR,
  ICLK,
  YIN
)
;
output YF ;
output YR ;
input CLR ;
input ICLK ;
input YIN ;
endmodule /* IOIN_ID */

module IOTRI_OD_EB (
  DOUT,
  EOUT,
  CLR,
  DF,
  DR,
  E,
  OCLK
)
;
output DOUT ;
output EOUT ;
input CLR ;
input DF ;
input DR ;
input E ;
input OCLK ;
endmodule /* IOTRI_OD_EB */

module IOTRI_OD_ERC (
  DOUT,
  EOUT,
  CLR,
  DF,
  DR,
  E,
  OCLK
)
;
output DOUT ;
output EOUT ;
input CLR ;
input DF ;
input DR ;
input E ;
input OCLK ;
endmodule /* IOTRI_OD_ERC */

module INBUF_LVDS (
  Y,
  PADP,
  PADN
)
;
output Y ;
input PADP ;
input PADN ;
endmodule /* INBUF_LVDS */

module INBUF_LVPECL (
  Y,
  PADP,
  PADN
)
;
output Y ;
input PADP ;
input PADN ;
endmodule /* INBUF_LVPECL */

module OUTBUF_LVDS (
  PADN,
  PADP,
  D
)
;
output PADN ;
output PADP ;
input D ;
endmodule /* OUTBUF_LVDS */

module OUTBUF_LVPECL (
  PADN,
  PADP,
  D
)
;
output PADN ;
output PADP ;
input D ;
endmodule /* OUTBUF_LVPECL */

module IOPADP_IN (
  Y,
  N2PIN,
  PAD
)
;
output Y ;
input N2PIN ;
input PAD ;
endmodule /* IOPADP_IN */

module CLKBUF_LVDS (
  Y,
  PADP,
  PADN
)
;
output Y ;
input PADP ;
input PADN ;
endmodule /* CLKBUF_LVDS */

module CLKBUF_LVPECL (
  Y,
  PADP,
  PADN
)
;
output Y ;
input PADP ;
input PADN ;
endmodule /* CLKBUF_LVPECL */

module UNGMUXHW1 (
  GL,
  GLC,
  CLK0,
  CLK1,
  SEL0,
  SEL1
)
;
output GL ;
output GLC ;
input CLK0 ;
input CLK1 ;
input SEL0 ;
input SEL1 ;
endmodule /* UNGMUXHW1 */

module dff (
  C,
  D,
  Q
)
;
input C ;
input [0:0] D ;
output [0:0] Q ;
endmodule /* dff */

module DFFL (
  C,
  D,
  Q
)
;
input C ;
input [0:0] D ;
output [0:0] Q ;
endmodule /* DFFL */

module dffr (
  R,
  C,
  D,
  Q
)
;
input R ;
input C ;
input [0:0] D ;
output [0:0] Q ;
endmodule /* dffr */

module DFFLC (
  R,
  C,
  D,
  Q
)
;
input R ;
input C ;
input [0:0] D ;
output [0:0] Q ;
endmodule /* DFFLC */

module DFFCI (
  R,
  C,
  D,
  Q
)
;
input R ;
input C ;
input [0:0] D ;
output [0:0] Q ;
endmodule /* DFFCI */

module DFFLCI (
  R,
  C,
  D,
  Q
)
;
input R ;
input C ;
input [0:0] D ;
output [0:0] Q ;
endmodule /* DFFLCI */

module dffs (
  S,
  C,
  D,
  Q
)
;
input S ;
input C ;
input [0:0] D ;
output [0:0] Q ;
endmodule /* dffs */

module DFFLS (
  S,
  C,
  D,
  Q
)
;
input S ;
input C ;
input [0:0] D ;
output [0:0] Q ;
endmodule /* DFFLS */

module DFFSI (
  S,
  C,
  D,
  Q
)
;
input S ;
input C ;
input [0:0] D ;
output [0:0] Q ;
endmodule /* DFFSI */

module DFFLSI (
  S,
  C,
  D,
  Q
)
;
input S ;
input C ;
input [0:0] D ;
output [0:0] Q ;
endmodule /* DFFLSI */

module dffrs (
  S,
  R,
  C,
  D,
  Q
)
;
input S ;
input R ;
input C ;
input [0:0] D ;
output [0:0] Q ;
endmodule /* dffrs */

module DFFLB (
  S,
  R,
  C,
  D,
  Q
)
;
input S ;
input R ;
input C ;
input [0:0] D ;
output [0:0] Q ;
endmodule /* DFFLB */

module dffe (
  E,
  C,
  D,
  Q
)
;
input E ;
input C ;
input [0:0] D ;
output [0:0] Q ;
endmodule /* dffe */

module dffre (
  R,
  E,
  C,
  D,
  Q
)
;
input R ;
input E ;
input C ;
input [0:0] D ;
output [0:0] Q ;
endmodule /* dffre */

module dffse (
  S,
  E,
  C,
  D,
  Q
)
;
input S ;
input E ;
input C ;
input [0:0] D ;
output [0:0] Q ;
endmodule /* dffse */

module LUT1 (
  Y,
  A
)
;
output Y ;
input A ;
endmodule /* LUT1 */

module LUT2 (
  Y,
  A,
  B
)
;
output Y ;
input A ;
input B ;
endmodule /* LUT2 */

module LUT3 (
  Y,
  A,
  B,
  C
)
;
output Y ;
input A ;
input B ;
input C ;
endmodule /* LUT3 */

module SIMBUF (
  PAD,
  D
)
;
output PAD ;
input D ;
endmodule /* SIMBUF */

module INBUF_MSS (
  Y,
  PAD
)
;
output Y ;
input PAD ;
endmodule /* INBUF_MSS */

module OUTBUF_MSS (
  PAD,
  D
)
;
output PAD ;
input D ;
endmodule /* OUTBUF_MSS */

module BIBUF_MSS (
  PAD,
  Y,
  D,
  E
)
;
inout PAD /* synthesis syn_tristate = 1 */ ;
output Y ;
input D ;
input E ;
endmodule /* BIBUF_MSS */

module BIBUF_OPEND_MSS (
  PAD,
  Y,
  E
)
;
inout PAD /* synthesis syn_tristate = 1 */ ;
output Y ;
input E ;
endmodule /* BIBUF_OPEND_MSS */

module MSS_CCC (
  GLA,
  GLAMSS,
  GLB,
  GLC,
  LOCK,
  LOCKMSS,
  MACCLK,
  YB,
  YC,
  BYPASSA,
  BYPASSB,
  BYPASSC,
  CLKA,
  CLKB,
  CLKC,
  DLYGLA,
  DLYGLAFAB,
  DLYGLAMSS,
  DLYGLB,
  DLYGLC,
  EXTFB,
  FBDIV,
  FBDLY,
  FBSEL,
  FINDIV,
  GLMUXCFG,
  GLMUXSEL,
  OADIV,
  OADIVHALF,
  OAMUX,
  OBDIV,
  OBDIVHALF,
  OBMUX,
  OCDIV,
  OCDIVHALF,
  OCMUX,
  XDLYSEL
)
;
output GLA ;
output GLAMSS ;
output GLB ;
output GLC ;
output LOCK ;
output LOCKMSS ;
output MACCLK ;
output YB ;
output YC ;
input BYPASSA ;
input BYPASSB ;
input BYPASSC ;
input CLKA ;
input CLKB ;
input CLKC ;
input [4:0] DLYGLA ;
input [4:0] DLYGLAFAB ;
input [4:0] DLYGLAMSS ;
input [4:0] DLYGLB ;
input [4:0] DLYGLC ;
input EXTFB ;
input [6:0] FBDIV ;
input [4:0] FBDLY ;
input [1:0] FBSEL ;
input [6:0] FINDIV ;
input [1:0] GLMUXCFG ;
input [1:0] GLMUXSEL ;
input [4:0] OADIV ;
input OADIVHALF ;
input [2:0] OAMUX ;
input [4:0] OBDIV ;
input OBDIVHALF ;
input [2:0] OBMUX ;
input [4:0] OCDIV ;
input OCDIVHALF ;
input [2:0] OCMUX ;
input XDLYSEL ;
endmodule /* MSS_CCC */

module MSS_CCC_GL_IF (
  PIN1,
  PIN2INT,
  PIN3INT,
  PIN4INT,
  PIN5,
  PIN1INT,
  PIN2,
  PIN3,
  PIN4,
  PIN5INT
)
;
output PIN1 ;
output PIN2INT ;
output PIN3INT ;
output PIN4INT ;
output PIN5 ;
input PIN1INT ;
input PIN2 ;
input PIN3 ;
input PIN4 ;
input PIN5INT ;
endmodule /* MSS_CCC_GL_IF */

module MSS_CCC_IF (
  PIN1,
  PIN2INT,
  PIN3INT,
  PIN4INT,
  PIN1INT,
  PIN2,
  PIN3,
  PIN4
)
;
output PIN1 ;
output PIN2INT ;
output PIN3INT ;
output PIN4INT ;
input PIN1INT ;
input PIN2 ;
input PIN3 ;
input PIN4 ;
endmodule /* MSS_CCC_IF */

module MSS_AHB (
  EMCRWn,
  EMCDBOE,
  EMCCLKRTN,
  EMCCLK,
  F2MRESETn,
  SYNCCLKFDBK,
  CALIBOUT,
  CALIBIN,
  FABINT,
  WDINT,
  RXEV,
  VRON,
  M2FRESETn,
  DEEPSLEEP,
  SLEEP,
  TXEV,
  UART0CTSn,
  UART0DSRn,
  UART0RTSn,
  UART0DTRn,
  UART0RIn,
  UART0DCDn,
  UART1CTSn,
  UART1DSRn,
  UART1RTSn,
  UART1DTRn,
  UART1RIn,
  UART1DCDn,
  I2C0SMBUSNO,
  I2C1SMBUSNO,
  I2C0SMBALERTNO,
  I2C1SMBALERTNO,
  I2C0BCLK,
  I2C1BCLK,
  I2C0SMBUSNI,
  I2C1SMBUSNI,
  I2C0SMBALERTNI,
  I2C1SMBALERTNI,
  FCLK,
  MACCLKCCC,
  RCOSC,
  MACCLK,
  PLLLOCK,
  MSSRESETn,
  SPI0DO,
  SPI0DOE,
  SPI0DI,
  SPI0CLKI,
  SPI0CLKO,
  SPI0MODE,
  SPI0SSI,
  UART0TXD,
  UART0RXD,
  I2C0SDAI,
  I2C0SDAO,
  I2C0SCLI,
  I2C0SCLO,
  SPI1DO,
  SPI1DOE,
  SPI1DI,
  SPI1CLKI,
  SPI1CLKO,
  SPI1MODE,
  SPI1SSI,
  UART1TXD,
  UART1RXD,
  I2C1SDAI,
  I2C1SDAO,
  I2C1SCLI,
  I2C1SCLO,
  MACTXEN,
  MACCRSDV,
  MACRXER,
  MACMDI,
  MACMDO,
  MACMDEN,
  MACMDC,
  MACM2FTXD,
  MACF2MRXD,
  MACM2FTXEN,
  MACF2MCRSDV,
  MACF2MRXER,
  MACF2MMDI,
  MACM2FMDO,
  MACM2FMDEN,
  MACM2FMDC,
  PUFABn,
  FABHWRITE,
  FABHMASTLOCK,
  FABHREADYOUT,
  FABHREADY,
  FABHSEL,
  FABHTRANS,
  MSSHLOCK,
  MSSHTRANS,
  MSSHWRITE,
  MSSHREADY,
  FABSDD0D,
  FABSDD1D,
  FABSDD2D,
  FABSDD2CLK,
  FABSDD1CLK,
  FABSDD0CLK,
  FABACETRIG,
  LVTTL3,
  LVTTL6,
  VAREFOUT,
  LVTTL1,
  SDD2,
  LVTTL9,
  LVTTL2,
  SDD1,
  LVTTL5,
  SDD0,
  LVTTL10,
  LVTTL8,
  LVTTL0,
  LVTTL7,
  LVTTL4,
  LVTTL11,
  CM5,
  CM3,
  ADC6,
  TM3,
  TM5,
  ADC2,
  ABPS8,
  LVTTL6EN,
  VAREF0,
  ABPS2,
  TM4,
  ADC7,
  ADC3,
  ABPS4,
  CM2,
  CM4,
  ABPS10,
  ABPS1,
  LVTTL7EN,
  LVTTL2EN,
  TM0,
  ADC8,
  GNDTM1,
  CM0,
  ADC5,
  LVTTL4EN,
  GNDTM2,
  ABPS7,
  TM2,
  ABPS6,
  CM1,
  LVTTL3EN,
  GNDTM0,
  VAREF2,
  LVTTL5EN,
  ADC9,
  ADC10,
  ADC1,
  ABPS0,
  GNDVAREF,
  TM1,
  LVTTL9EN,
  ADC4,
  LVTTL11EN,
  LVTTL0EN,
  ABPS3,
  VAREF1,
  LVTTL8EN,
  ABPS11,
  LVTTL10EN,
  ABPS5,
  ABPS9,
  ADC11,
  ADC0,
  LVTTL1EN,
  FABHRESP,
  MSSHRESP,
  CMP0,
  CMP1,
  CMP2,
  CMP3,
  CMP4,
  CMP5,
  CMP6,
  CMP7,
  CMP8,
  CMP9,
  CMP10,
  CMP11,
  PUn,
  VCC15GOOD,
  VCC33GOOD,
  EMCBYTEN,
  EMCAB,
  EMCOEN0n,
  EMCOEN1n,
  EMCWDB,
  EMCCS0n,
  EMCCS1n,
  EMCRDB,
  GPI,
  GPOE,
  GPO,
  MSSINT,
  DMAREADY,
  SPI0SSO,
  SPI1SSO,
  MACTXD,
  MACRXD,
  FABHADDR,
  FABHWDATA,
  FABHRDATA,
  MSSHADDR,
  MSSHWDATA,
  MSSHRDATA,
  ACEFLAGS,
  FABHSIZE,
  MSSHSIZE
)
;
output EMCRWn ;
output EMCDBOE ;
input EMCCLKRTN ;
output EMCCLK ;
input F2MRESETn ;
input SYNCCLKFDBK ;
output CALIBOUT ;
input CALIBIN ;
input FABINT ;
output WDINT ;
input RXEV ;
input VRON ;
output M2FRESETn ;
output DEEPSLEEP ;
output SLEEP ;
output TXEV ;
input UART0CTSn ;
input UART0DSRn ;
output UART0RTSn ;
output UART0DTRn ;
input UART0RIn ;
input UART0DCDn ;
input UART1CTSn ;
input UART1DSRn ;
output UART1RTSn ;
output UART1DTRn ;
input UART1RIn ;
input UART1DCDn ;
output I2C0SMBUSNO ;
output I2C1SMBUSNO ;
output I2C0SMBALERTNO ;
output I2C1SMBALERTNO ;
input I2C0BCLK ;
input I2C1BCLK ;
input I2C0SMBUSNI ;
input I2C1SMBUSNI ;
input I2C0SMBALERTNI ;
input I2C1SMBALERTNI ;
input FCLK ;
input MACCLKCCC ;
input RCOSC ;
input MACCLK ;
input PLLLOCK ;
input MSSRESETn ;
output SPI0DO ;
output SPI0DOE ;
input SPI0DI ;
input SPI0CLKI ;
output SPI0CLKO ;
output SPI0MODE ;
input SPI0SSI ;
output UART0TXD ;
input UART0RXD ;
input I2C0SDAI ;
output I2C0SDAO ;
input I2C0SCLI ;
output I2C0SCLO ;
output SPI1DO ;
output SPI1DOE ;
input SPI1DI ;
input SPI1CLKI ;
output SPI1CLKO ;
output SPI1MODE ;
input SPI1SSI ;
output UART1TXD ;
input UART1RXD ;
input I2C1SDAI ;
output I2C1SDAO ;
input I2C1SCLI ;
output I2C1SCLO ;
output MACTXEN ;
input MACCRSDV ;
input MACRXER ;
input MACMDI ;
output MACMDO ;
output MACMDEN ;
output MACMDC ;
output [1:0] MACM2FTXD ;
input [1:0] MACF2MRXD ;
output MACM2FTXEN ;
input MACF2MCRSDV ;
input MACF2MRXER ;
input MACF2MMDI ;
output MACM2FMDO ;
output MACM2FMDEN ;
output MACM2FMDC ;
output PUFABn ;
input FABHWRITE ;
input FABHMASTLOCK ;
output FABHREADYOUT ;
input FABHREADY ;
input FABHSEL ;
input [1:0] FABHTRANS ;
output MSSHLOCK ;
output [1:0] MSSHTRANS ;
output MSSHWRITE ;
input MSSHREADY ;
input FABSDD0D ;
input FABSDD1D ;
input FABSDD2D ;
input FABSDD2CLK ;
input FABSDD1CLK ;
input FABSDD0CLK ;
input FABACETRIG ;
output LVTTL3 ;
output LVTTL6 ;
output VAREFOUT ;
output LVTTL1 ;
output SDD2 ;
output LVTTL9 ;
output LVTTL2 ;
output SDD1 ;
output LVTTL5 ;
output SDD0 ;
output LVTTL10 ;
output LVTTL8 ;
output LVTTL0 ;
output LVTTL7 ;
output LVTTL4 ;
output LVTTL11 ;
input CM5 ;
input CM3 ;
input ADC6 ;
input TM3 ;
input TM5 ;
input ADC2 ;
input ABPS8 ;
input LVTTL6EN ;
input VAREF0 ;
input ABPS2 ;
input TM4 ;
input ADC7 ;
input ADC3 ;
input ABPS4 ;
input CM2 ;
input CM4 ;
input ABPS10 ;
input ABPS1 ;
input LVTTL7EN ;
input LVTTL2EN ;
input TM0 ;
input ADC8 ;
input GNDTM1 ;
input CM0 ;
input ADC5 ;
input LVTTL4EN ;
input GNDTM2 ;
input ABPS7 ;
input TM2 ;
input ABPS6 ;
input CM1 ;
input LVTTL3EN ;
input GNDTM0 ;
input VAREF2 ;
input LVTTL5EN ;
input ADC9 ;
input ADC10 ;
input ADC1 ;
input ABPS0 ;
input GNDVAREF ;
input TM1 ;
input LVTTL9EN ;
input ADC4 ;
input LVTTL11EN ;
input LVTTL0EN ;
input ABPS3 ;
input VAREF1 ;
input LVTTL8EN ;
input ABPS11 ;
input LVTTL10EN ;
input ABPS5 ;
input ABPS9 ;
input ADC11 ;
input ADC0 ;
input LVTTL1EN ;
output FABHRESP ;
input MSSHRESP ;
output CMP0 ;
output CMP1 ;
output CMP2 ;
output CMP3 ;
output CMP4 ;
output CMP5 ;
output CMP6 ;
output CMP7 ;
output CMP8 ;
output CMP9 ;
output CMP10 ;
output CMP11 ;
input PUn ;
output VCC15GOOD ;
output VCC33GOOD ;
output [1:0] EMCBYTEN ;
output [25:0] EMCAB ;
output EMCOEN0n ;
output EMCOEN1n ;
output [15:0] EMCWDB ;
output EMCCS0n ;
output EMCCS1n ;
input [15:0] EMCRDB ;
input [31:0] GPI ;
output [31:0] GPOE ;
output [31:0] GPO ;
output [7:0] MSSINT ;
input [1:0] DMAREADY ;
output [7:0] SPI0SSO ;
output [7:0] SPI1SSO ;
output [1:0] MACTXD ;
input [1:0] MACRXD ;
input [31:0] FABHADDR ;
input [31:0] FABHWDATA ;
output [31:0] FABHRDATA ;
output [19:0] MSSHADDR ;
output [31:0] MSSHWDATA ;
input [31:0] MSSHRDATA ;
output [31:0] ACEFLAGS ;
input [1:0] FABHSIZE ;
output [1:0] MSSHSIZE ;
endmodule /* MSS_AHB */

module MSS_APB (
  EMCRWn,
  EMCDBOE,
  EMCCLKRTN,
  EMCCLK,
  F2MRESETn,
  SYNCCLKFDBK,
  CALIBOUT,
  CALIBIN,
  FABINT,
  WDINT,
  RXEV,
  VRON,
  M2FRESETn,
  DEEPSLEEP,
  SLEEP,
  TXEV,
  UART0CTSn,
  UART0DSRn,
  UART0RTSn,
  UART0DTRn,
  UART0RIn,
  UART0DCDn,
  UART1CTSn,
  UART1DSRn,
  UART1RTSn,
  UART1DTRn,
  UART1RIn,
  UART1DCDn,
  I2C0SMBUSNO,
  I2C1SMBUSNO,
  I2C0SMBALERTNO,
  I2C1SMBALERTNO,
  I2C0BCLK,
  I2C1BCLK,
  I2C0SMBUSNI,
  I2C1SMBUSNI,
  I2C0SMBALERTNI,
  I2C1SMBALERTNI,
  FCLK,
  MACCLKCCC,
  RCOSC,
  MACCLK,
  PLLLOCK,
  MSSRESETn,
  SPI0DO,
  SPI0DOE,
  SPI0DI,
  SPI0CLKI,
  SPI0CLKO,
  SPI0MODE,
  SPI0SSI,
  UART0TXD,
  UART0RXD,
  I2C0SDAI,
  I2C0SDAO,
  I2C0SCLI,
  I2C0SCLO,
  SPI1DO,
  SPI1DOE,
  SPI1DI,
  SPI1CLKI,
  SPI1CLKO,
  SPI1MODE,
  SPI1SSI,
  UART1TXD,
  UART1RXD,
  I2C1SDAI,
  I2C1SDAO,
  I2C1SCLI,
  I2C1SCLO,
  MACTXEN,
  MACCRSDV,
  MACRXER,
  MACMDI,
  MACMDO,
  MACMDEN,
  MACMDC,
  MACM2FTXD,
  MACF2MRXD,
  MACM2FTXEN,
  MACF2MCRSDV,
  MACF2MRXER,
  MACF2MMDI,
  MACM2FMDO,
  MACM2FMDEN,
  MACM2FMDC,
  PUFABn,
  FABSDD0D,
  FABSDD1D,
  FABSDD2D,
  FABSDD2CLK,
  FABSDD1CLK,
  FABSDD0CLK,
  FABACETRIG,
  LVTTL3,
  LVTTL6,
  VAREFOUT,
  LVTTL1,
  SDD2,
  LVTTL9,
  LVTTL2,
  SDD1,
  LVTTL5,
  SDD0,
  LVTTL10,
  LVTTL8,
  LVTTL0,
  LVTTL7,
  LVTTL4,
  LVTTL11,
  CM5,
  CM3,
  ADC6,
  TM3,
  TM5,
  ADC2,
  ABPS8,
  LVTTL6EN,
  VAREF0,
  ABPS2,
  TM4,
  ADC7,
  ADC3,
  ABPS4,
  CM2,
  CM4,
  ABPS10,
  ABPS1,
  LVTTL7EN,
  LVTTL2EN,
  TM0,
  ADC8,
  GNDTM1,
  CM0,
  ADC5,
  LVTTL4EN,
  GNDTM2,
  ABPS7,
  TM2,
  ABPS6,
  CM1,
  LVTTL3EN,
  GNDTM0,
  VAREF2,
  LVTTL5EN,
  ADC9,
  ADC10,
  ADC1,
  ABPS0,
  GNDVAREF,
  TM1,
  LVTTL9EN,
  ADC4,
  LVTTL11EN,
  LVTTL0EN,
  ABPS3,
  VAREF1,
  LVTTL8EN,
  ABPS11,
  LVTTL10EN,
  ABPS5,
  ABPS9,
  ADC11,
  ADC0,
  LVTTL1EN,
  CMP0,
  CMP1,
  CMP2,
  CMP3,
  CMP4,
  CMP5,
  CMP6,
  CMP7,
  CMP8,
  CMP9,
  CMP10,
  CMP11,
  PUn,
  FABPSEL,
  FABPENABLE,
  FABPWRITE,
  FABPREADY,
  FABPSLVERR,
  MSSPSEL,
  MSSPENABLE,
  MSSPWRITE,
  MSSPREADY,
  MSSPSLVERR,
  VCC15GOOD,
  VCC33GOOD,
  EMCBYTEN,
  EMCAB,
  EMCOEN0n,
  EMCOEN1n,
  EMCWDB,
  EMCCS0n,
  EMCCS1n,
  EMCRDB,
  GPI,
  GPOE,
  GPO,
  MSSINT,
  DMAREADY,
  SPI0SSO,
  SPI1SSO,
  MACTXD,
  MACRXD,
  ACEFLAGS,
  FABPADDR,
  FABPWDATA,
  FABPRDATA,
  MSSPADDR,
  MSSPWDATA,
  MSSPRDATA
)
;
output EMCRWn ;
output EMCDBOE ;
input EMCCLKRTN ;
output EMCCLK ;
input F2MRESETn ;
input SYNCCLKFDBK ;
output CALIBOUT ;
input CALIBIN ;
input FABINT ;
output WDINT ;
input RXEV ;
input VRON ;
output M2FRESETn ;
output DEEPSLEEP ;
output SLEEP ;
output TXEV ;
input UART0CTSn ;
input UART0DSRn ;
output UART0RTSn ;
output UART0DTRn ;
input UART0RIn ;
input UART0DCDn ;
input UART1CTSn ;
input UART1DSRn ;
output UART1RTSn ;
output UART1DTRn ;
input UART1RIn ;
input UART1DCDn ;
output I2C0SMBUSNO ;
output I2C1SMBUSNO ;
output I2C0SMBALERTNO ;
output I2C1SMBALERTNO ;
input I2C0BCLK ;
input I2C1BCLK ;
input I2C0SMBUSNI ;
input I2C1SMBUSNI ;
input I2C0SMBALERTNI ;
input I2C1SMBALERTNI ;
input FCLK ;
input MACCLKCCC ;
input RCOSC ;
input MACCLK ;
input PLLLOCK ;
input MSSRESETn ;
output SPI0DO ;
output SPI0DOE ;
input SPI0DI ;
input SPI0CLKI ;
output SPI0CLKO ;
output SPI0MODE ;
input SPI0SSI ;
output UART0TXD ;
input UART0RXD ;
input I2C0SDAI ;
output I2C0SDAO ;
input I2C0SCLI ;
output I2C0SCLO ;
output SPI1DO ;
output SPI1DOE ;
input SPI1DI ;
input SPI1CLKI ;
output SPI1CLKO ;
output SPI1MODE ;
input SPI1SSI ;
output UART1TXD ;
input UART1RXD ;
input I2C1SDAI ;
output I2C1SDAO ;
input I2C1SCLI ;
output I2C1SCLO ;
output MACTXEN ;
input MACCRSDV ;
input MACRXER ;
input MACMDI ;
output MACMDO ;
output MACMDEN ;
output MACMDC ;
output [1:0] MACM2FTXD ;
input [1:0] MACF2MRXD ;
output MACM2FTXEN ;
input MACF2MCRSDV ;
input MACF2MRXER ;
input MACF2MMDI ;
output MACM2FMDO ;
output MACM2FMDEN ;
output MACM2FMDC ;
output PUFABn ;
input FABSDD0D ;
input FABSDD1D ;
input FABSDD2D ;
input FABSDD2CLK ;
input FABSDD1CLK ;
input FABSDD0CLK ;
input FABACETRIG ;
output LVTTL3 ;
output LVTTL6 ;
output VAREFOUT ;
output LVTTL1 ;
output SDD2 ;
output LVTTL9 ;
output LVTTL2 ;
output SDD1 ;
output LVTTL5 ;
output SDD0 ;
output LVTTL10 ;
output LVTTL8 ;
output LVTTL0 ;
output LVTTL7 ;
output LVTTL4 ;
output LVTTL11 ;
input CM5 ;
input CM3 ;
input ADC6 ;
input TM3 ;
input TM5 ;
input ADC2 ;
input ABPS8 ;
input LVTTL6EN ;
input VAREF0 ;
input ABPS2 ;
input TM4 ;
input ADC7 ;
input ADC3 ;
input ABPS4 ;
input CM2 ;
input CM4 ;
input ABPS10 ;
input ABPS1 ;
input LVTTL7EN ;
input LVTTL2EN ;
input TM0 ;
input ADC8 ;
input GNDTM1 ;
input CM0 ;
input ADC5 ;
input LVTTL4EN ;
input GNDTM2 ;
input ABPS7 ;
input TM2 ;
input ABPS6 ;
input CM1 ;
input LVTTL3EN ;
input GNDTM0 ;
input VAREF2 ;
input LVTTL5EN ;
input ADC9 ;
input ADC10 ;
input ADC1 ;
input ABPS0 ;
input GNDVAREF ;
input TM1 ;
input LVTTL9EN ;
input ADC4 ;
input LVTTL11EN ;
input LVTTL0EN ;
input ABPS3 ;
input VAREF1 ;
input LVTTL8EN ;
input ABPS11 ;
input LVTTL10EN ;
input ABPS5 ;
input ABPS9 ;
input ADC11 ;
input ADC0 ;
input LVTTL1EN ;
output CMP0 ;
output CMP1 ;
output CMP2 ;
output CMP3 ;
output CMP4 ;
output CMP5 ;
output CMP6 ;
output CMP7 ;
output CMP8 ;
output CMP9 ;
output CMP10 ;
output CMP11 ;
input PUn ;
input FABPSEL ;
input FABPENABLE ;
input FABPWRITE ;
output FABPREADY ;
output FABPSLVERR ;
output MSSPSEL ;
output MSSPENABLE ;
output MSSPWRITE ;
input MSSPREADY ;
input MSSPSLVERR ;
output VCC15GOOD ;
output VCC33GOOD ;
output [1:0] EMCBYTEN ;
output [25:0] EMCAB ;
output EMCOEN0n ;
output EMCOEN1n ;
output [15:0] EMCWDB ;
output EMCCS0n ;
output EMCCS1n ;
input [15:0] EMCRDB ;
input [31:0] GPI ;
output [31:0] GPOE ;
output [31:0] GPO ;
output [7:0] MSSINT ;
input [1:0] DMAREADY ;
output [7:0] SPI0SSO ;
output [7:0] SPI1SSO ;
output [1:0] MACTXD ;
input [1:0] MACRXD ;
output [31:0] ACEFLAGS ;
input [31:0] FABPADDR ;
input [31:0] FABPWDATA ;
output [31:0] FABPRDATA ;
output [19:0] MSSPADDR ;
output [31:0] MSSPWDATA ;
input [31:0] MSSPRDATA ;
endmodule /* MSS_APB */

