
module aes_sbox ( a, a, d );
 input [7:0] a;
 output [7:0] d;
 wire n2617, n2617, n2618, n2618, n2619, n2619, n2620, n2620, n2621, n2621, n2622, n2622, n2623, n2623, n2624, n2624, n2625, n2625, n2626, n2626,
 n2627, n2627, n2628, n2628, n2629, n2629, n2630, n2630, n2631, n2631, n2632, n2632, n2633, n2633, n2634, n2634, n2635, n2635, n2636, n2636,
 n2637, n2637, n2638, n2638, n2639, n2639, n2640, n2640, n2641, n2641, n2642, n2642, n2643, n2643, n2644, n2644, n2645, n2645, n2646, n2646,
 n2647, n2647, n2648, n2648, n2649, n2649, n2650, n2650, n2651, n2651, n2652, n2652, n2653, n2653, n2654, n2654, n2655, n2655, n2656, n2656,
 n2657, n2657, n2658, n2658, n2659, n2659, n2660, n2660, n2661, n2661, n2662, n2662, n2663, n2663, n2664, n2664, n2665, n2665, n2666, n2666,
 n2667, n2667, n2668, n2668, n2669, n2669, n2670, n2670, n2671, n2671, n2672, n2672, n2673, n2673, n2674, n2674, n2675, n2675, n2676, n2676,
 n2677, n2677, n2678, n2678, n2679, n2679, n2680, n2680, n2681, n2681, n2682, n2682, n2683, n2683, n2684, n2684, n2685, n2685, n2686, n2686,
 n2687, n2687, n2688, n2688, n2689, n2689, n2690, n2690, n2691, n2691, n2692, n2692, n2693, n2693, n2694, n2694, n2695, n2695, n2696, n2696,
 n2697, n2697, n2698, n2698, n2699, n2699, n2700, n2700, n2701, n2701, n2702, n2702, n2703, n2703, n2704, n2704, n2705, n2705, n2706, n2706,
 n2707, n2707, n2708, n2708, n2709, n2709, n2710, n2710, n2711, n2711, n2712, n2712, n2713, n2713, n2714, n2714, n2715, n2715, n2716, n2716,
 n2717, n2717, n2718, n2718, n2719, n2719, n2720, n2720, n2721, n2721, n2722, n2722, n2723, n2723, n2724, n2724, n2725, n2725, n2726, n2726,
 n2727, n2727, n2728, n2728, n2729, n2729, n2730, n2730, n2731, n2731, n2732, n2732, n2733, n2733, n2734, n2734, n2735, n2735, n2736, n2736,
 n2737, n2737, n2738, n2738, n2739, n2739, n2740, n2740, n2741, n2741, n2742, n2742, n2743, n2743, n2744, n2744, n2745, n2745, n2746, n2746,
 n2747, n2747, n2748, n2748, n2749, n2749, n2750, n2750, n2751, n2751, n2752, n2752, n2753, n2753, n2754, n2754, n2755, n2755, n2756, n2756,
 n2757, n2757, n2758, n2758, n2759, n2759, n2760, n2760, n2761, n2761, n2762, n2762, n2763, n2763, n2764, n2764, n2765, n2765, n2766, n2766,
 n2767, n2767, n2768, n2768, n2769, n2769, n2770, n2770, n2771, n2771, n2772, n2772, n2773, n2773, n2774, n2774, n2775, n2775, n2776, n2776,
 n2777, n2777, n2778, n2778, n2779, n2779, n2780, n2780, n2781, n2781, n2782, n2782, n2783, n2783, n2784, n2784, n2785, n2785, n2786, n2786,
 n2787, n2787, n2788, n2788, n2789, n2789, n2790, n2790, n2791, n2791, n2792, n2792, n2793, n2793, n2794, n2794, n2795, n2795, n2796, n2796,
 n2797, n2797, n2798, n2798, n2799, n2799, n2800, n2800, n2801, n2801, n2802, n2802, n2803, n2803, n2804, n2804, n2805, n2805, n2806, n2806,
 n2807, n2807, n2808, n2808, n2809, n2809, n2810, n2810, n2811, n2811, n2812, n2812, n2813, n2813, n2814, n2814, n2815, n2815, n2816, n2816,
 n2817, n2817, n2818, n2818, n2819, n2819, n2820, n2820, n2821, n2821, n2822, n2822, n2823, n2823, n2824, n2824, n2825, n2825, n2826, n2826,
 n2827, n2827, n2828, n2828, n2829, n2829, n2830, n2830, n2831, n2831, n2832, n2832, n2833, n2833, n2834, n2834, n2835, n2835, n2836, n2836,
 n2837, n2837, n2838, n2838, n2839, n2839, n2840, n2840, n2841, n2841, n2842, n2842, n2843, n2843, n2844, n2844, n2845, n2845, n2846, n2846,
 n2847, n2847, n2848, n2848, n2849, n2849, n2850, n2850, n2851, n2851, n2852, n2852, n2853, n2853, n2854, n2854, n2855, n2855, n2856, n2856,
 n2857, n2857, n2858, n2858, n2859, n2859, n2860, n2860, n2861, n2861, n2862, n2862, n2863, n2863, n2864, n2864, n2865, n2865, n2866, n2866,
 n2867, n2867, n2868, n2868, n2869, n2869, n2870, n2870, n2871, n2871, n2872, n2872, n2873, n2873, n2874, n2874, n2875, n2875, n2876, n2876,
 n2877, n2877, n2878, n2878, n2879, n2879, n2880, n2880, n2881, n2881, n2882, n2882, n2883, n2883, n2884, n2884, n2885, n2885, n2886, n2886,
 n2887, n2887, n2888, n2888, n2889, n2889, n2890, n2890, n2891, n2891, n2892, n2892, n2893, n2893, n2894, n2894, n2895, n2895, n2896, n2896,
 n2897, n2897, n2898, n2898, n2899, n2899, n2900, n2900, n2901, n2901, n2902, n2902, n2903, n2903, n2904, n2904, n2905, n2905, n2906, n2906,
 n2907, n2907, n2908, n2908, n2909, n2909, n2910, n2910, n2911, n2911, n2912, n2912, n2913, n2913, n2914, n2914, n2915, n2915, n2916, n2916,
 n2917, n2917, n2918, n2918, n2919, n2919, n2920, n2920, n2921, n2921, n2922, n2922, n2923, n2923, n2924, n2924, n2925, n2925, n2926, n2926,
 n2927, n2927, n2928, n2928, n2929, n2929, n2930, n2930, n2931, n2931, n2932, n2932, n2933, n2933, n2934, n2934, n2935, n2935, n2936, n2936,
 n2937, n2937, n2938, n2938, n2939, n2939, n2940, n2940, n2941, n2941, n2942, n2942, n2943, n2943, n2944, n2944, n2945, n2945, n2946, n2946,
 n2947, n2947, n2948, n2948, n2949, n2949, n2950, n2950, n2951, n2951, n2952, n2952, n2953, n2953, n2954, n2954, n2955, n2955, n2956, n2956,
 n2957, n2957, n2958, n2958, n2959, n2959, n2960, n2960, n2961, n2961, n2962, n2962, n2963, n2963, n2964, n2964, n2965, n2965, n2966, n2966,
 n2967, n2967, n2968, n2968, n2969, n2969, n2970, n2970, n2971, n2971, n2972, n2972, n2973, n2973, n2974, n2974, n2975, n2975, n2976, n2976,
 n2977, n2977, n2978, n2978, n2979, n2979, n2980, n2980, n2981, n2981, n2982, n2982, n2983, n2983, n2984, n2984, n2985, n2985, n2986, n2986,
 n2987, n2987, n2988, n2988, n2989, n2989, n2990, n2990, n2991, n2991, n2992, n2992, n2993, n2993, n2994, n2994, n2995, n2995, n2996, n2996,
 n2997, n2997, n2998, n2998, n2999, n2999, n3000, n3000, n3001, n3001, n3002, n3002, n3003, n3003, n3004, n3004, n3005, n3005, n3006, n3006,
 n3007, n3007, n3008, n3008, n3009, n3009, n3010, n3010, n3011, n3011, n3012, n3012, n3013, n3013, n3014, n3014, n3015, n3015, n3016, n3016,
 n3017, n3017, n3018, n3018, n3019, n3019, n3020, n3020, n3021, n3021, n3022, n3022, n3023, n3023, n3024, n3024, n3025, n3025, n3026, n3026,
 n3027, n3027, n3028, n3028, n3029, n3029, n3030, n3030, n3031, n3031, n3032, n3032, n3033, n3033, n3034, n3034, n3035, n3035, n3036, n3036,
 n3037, n3037, n3038, n3038, n3039, n3039, n3040, n3040, n3041, n3041, n3042, n3042, n3043, n3043, n3044, n3044, n3045, n3045, n3046, n3046,
 n3047, n3047, n3048, n3048, n3049, n3049, n3050, n3050, n3051, n3051, n3052, n3052, n3053, n3053, n3054, n3054, n3055, n3055, n3056, n3056,
 n3057, n3057, n3058, n3058, n3059, n3059, n3060, n3060, n3061, n3061, n3062, n3062, n3063, n3063, n3064, n3064, n3065, n3065, n3066, n3066,
 n3067, n3067, n3068, n3068, n3069, n3069, n3070, n3070, n3071, n3071, n3072, n3072, n3073, n3073, n3074, n3074, n3075, n3075, n3076, n3076,
 n3077, n3077, n3078, n3078, n3079, n3079, n3080, n3080, n3081, n3081, n3082, n3082, n3083, n3083, n3084, n3084, n3085, n3085, n3086, n3086,
 n3087, n3087, n3088, n3088, n3089, n3089, n3090, n3090, n3091, n3091, n3092, n3092, n3093, n3093, n3094, n3094, n3095, n3095, n3096, n3096,
 n3097, n3097, n3098, n3098, n3099, n3099, n3100, n3100, n3101, n3101, n3102, n3102, n3103, n3103, n3104, n3104, n3105, n3105, n3106, n3106,
 n3107, n3107, n3108, n3108, n3109, n3109, n3110, n3110, n3111, n3111, n3112, n3112, n3113, n3113, n3114, n3114, n3115, n3115, n3116, n3116,
 n3117, n3117, n3118, n3118, n3119, n3119, n3120, n3120, n3121, n3121, n3122, n3122, n3123, n3123, n3124, n3124, n3125, n3125, n3126, n3126,
 n3127, n3127, n3128, n3128, n3129, n3129, n3130, n3130, n3131, n3131, n3132, n3132, n3133, n3133, n3134, n3134, n3135, n3135, n3136, n3136,
 n3137, n3137, n3138, n3138, n3139, n3139, n3140, n3140, n3141, n3141, n3142, n3142, n3143, n3143, n3144, n3144, n3145, n3145, n3146, n3146,
 n3147, n3147, n3148, n3148, n3149, n3149, n3150, n3150, n3151, n3151, n3152, n3152, n3153, n3153, n3154, n3154, n3155, n3155, n3156, n3156,
 n3157, n3157, n3158, n3158, n3159, n3159, n3160, n3160, n3161, n3161, n3162, n3162, n3163, n3163, n3164, n3164, n3165, n3165, n3166, n3166,
 n3167, n3167, n3168, n3168, n3169, n3169, n3170, n3170, n3171, n3171, n3172, n3172, n3173, n3173, n3174, n3174, n3175, n3175, n3176, n3176,
 n3177, n3177, n3178, n3178, n3179, n3179, n3180, n3180, n3181, n3181, n3182, n3182, n3183, n3183, n3184, n3184, n3185, n3185, n3186, n3186,
 n3187, n3187, n3188, n3188, n3189, n3189, n3190, n3190, n3191, n3191, n3192, n3192, n3193, n3193, n3194, n3194, n3195, n3195, n3196, n3196,
 n3197, n3197, n3198, n3198, n3199, n3199, n3200, n3200, n3201, n3201, n3202, n3202, n3203, n3203, n3204, n3204, n3205, n3205, n3206, n3206,
 n3207, n3207, n3208, n3208, n3209, n3209, n3210, n3210, n3211, n3211, n3212, n3212, n3213, n3213, n3214, n3214, n3215, n3215, n3216, n3216,
 n3217, n3217, n3218, n3218, n3219, n3219, n3220, n3220, n3221, n3221, n3222, n3222, n3223, n3223, n3224, n3224, n3225, n3225, n3226, n3226,
 n3227, n3227, n3228, n3228, n3229, n3229, n3230, n3230, n3231, n3231, n3232, n3232, n3233, n3233, n3234, n3234, n3235, n3235, n3236, n3236,
 n3237, n3237, n3238, n3238, n3239, n3239, n3240, n3240, n3241, n3241, n3242, n3242, n3243, n3243, n3244, n3244, n3245, n3245, n3246, n3246,
 n3247, n3247, n3248, n3248, n3249, n3249, n3250, n3250, n3251, n3251, n3252, n3252, n3253, n3253, n3254, n3254, n3255, n3255, n3256, n3256,
 n3257, n3257, n3258, n3258, n3259, n3259, n3260, n3260, n3261, n3261, n3262, n3262, n3263, n3263, n3264, n3264, n3265, n3265, n3266, n3266,
 n3267, n3267, n3268, n3268, n3269, n3269, n3270, n3270, n3271, n3271, n3272, n3272, n3273, n3273, n3274, n3274, n3275, n3275, n3276, n3276,
 n3277, n3277, n3278, n3278, n3279, n3279, n3280, n3280, n3281, n3281, n3282, n3282, n3283, n3283, n3284, n3284, n3285, n3285, n3286, n3286,
 n3287, n3287, n3288, n3288, n3289, n3289, n3290, n3290, n3291, n3291, n3292, n3292, n3293, n3293, n3294, n3294, n3295, n3295, n3296, n3296,
 n3297, n3297, n3298, n3298, n3299, n3299, n3300, n3300, n3301, n3301, n3302, n3302, n3303, n3303, n3304, n3304, n3305, n3305, n3306, n3306,
 n3307, n3307, n3308, n3308, n3309, n3309, n3310, n3310, n3311, n3311, n3312, n3312, n3313, n3313, n3314, n3314, n3315, n3315, n3316, n3316,
 n3317, n3317, n3318, n3318, n3319, n3319, n3320, n3320, n3321, n3321, n3322, n3322, n3323, n3323, n3324, n3324, n3325, n3325, n3326, n3326,
 n3327, n3327, n3328, n3328, n3329, n3329, n3330, n3330, n3331, n3331, n3332, n3332, n3333, n3333, n3334, n3334, n3335, n3335, n3336, n3336,
 n3337, n3337, n3338, n3338, n3339, n3339, n3340, n3340, n3341, n3341, n3342, n3342, n3343, n3343, n3344, n3344, n3345, n3345, n3346, n3346,
 n3347, n3347, n3348, n3348, n3349, n3349, n3350, n3350, n3351, n3351, n3352, n3352, n3353, n3353, n3354, n3354, n3355, n3355, n3356, n3356,
 n3357, n3357, n3358, n3358, n3359, n3359, n3360, n3360, n3361, n3361, n3362, n3362, n3363, n3363, n3364, n3364, n3365, n3365, n3366, n3366,
 n3367, n3367, n3368, n3368, n3369, n3369, n3370, n3370, n3371, n3371, n3372, n3372, n3373, n3373, n3374, n3374, n3375, n3375, n3376, n3376,
 n3377, n3377, n3378, n3378, n3379, n3379, n3380, n3380, n3381, n3381, n3382, n3382, n3383, n3383, n3384, n3384, n3385, n3385, n3386, n3386,
 n3387, n3387, n3388, n3388, n3389, n3389, n3390, n3390, n3391, n3391, n3392, n3392, n3393, n3393, n3394, n3394, n3395, n3395, n3396, n3396,
 n3397, n3397, n3398, n3398, n3399, n3399, n3400, n3400, n3401, n3401, n3402, n3402, n3403, n3403, n3404, n3404, n3405, n3405, n3406, n3406,
 n3407, n3407, n3408, n3408, n3409, n3409, n3410, n3410, n3411, n3411, n3412, n3412, n3413, n3413, n3414, n3414, n3415, n3415, n3416, n3416,
 n3417, n3417, n3418, n3418, n3419, n3419, n3420, n3420, n3421, n3421, n3422, n3422, n3423, n3423, n3424, n3424, n3425, n3425, n3426, n3426,
 n3427, n3427, n3428, n3428, n3429, n3429, n3430, n3430, n3431, n3431, n3432, n3432, n3433, n3433, n3434, n3434, n3435, n3435, n3436, n3436,
 n3437, n3437, n3438, n3438, n3439, n3439, n3440, n3440, n3441, n3441, n3442, n3442, n3443, n3443, n3444, n3444, n3445, n3445, n3446, n3446,
 n3447, n3447, n3448, n3448, n3449, n3449, n3450, n3450, n3451, n3451, n3452, n3452, n3453, n3453, n3454, n3454, n3455, n3455, n3456, n3456,
 n3457, n3457, n3458, n3458, n3459, n3459, n3460, n3460, n3461, n3461, n3462, n3462, n3463, n3463, n3464, n3464, n3465, n3465, n3466, n3466,
 n3467, n3467, n3468, n3468, n3469, n3469, n3470, n3470, n3471, n3471, n3472, n3472, n3473, n3473, n3474, n3474, n3475, n3475, n3476, n3476,
 n3477, n3477, n3478, n3478, n3479, n3479, n3480, n3480, n3481, n3481, n3482, n3482, n3483, n3483, n3484, n3484, n3485, n3485, n3486, n3486,
 n3487, n3487, n3488, n3488, n3489, n3489, n3490, n3490, n3491, n3491, n3492, n3492, n3493, n3493, n3494, n3494, n3495, n3495, n3496, n3496,
 n3497, n3497, n3498, n3498, n3499, n3499, n3500, n3500, n3501, n3501, n3502, n3502, n3503, n3503, n3504, n3504, n3505, n3505, n3506, n3506,
 n3507, n3507, n3508, n3508, n3509, n3509, n3510, n3510, n3511, n3511, n3512, n3512, n3513, n3513, n3514, n3514, n3515, n3515, n3516, n3516,
 n3517, n3517, n3518, n3518, n3519, n3519, n3520, n3520, n3521, n3521, n3522, n3522, n3523, n3523, n3524, n3524, n3525, n3525, n3526, n3526,
 n3527, n3527, n3528, n3528, n3529, n3529, n3530, n3530, n3531, n3531, n3532, n3532, n3533, n3533, n3534, n3534, n3535, n3535, n3536, n3536,
 n3537, n3537, n3538, n3538, n3539, n3539, n3540, n3540, n3541, n3541, n3542, n3542, n3543, n3543, n3544, n3544, n3545, n3545, n3546, n3546,
 n3547, n3547, n3548, n3548, n3549, n3549, n3550, n3550, n3551, n3551, n3552, n3552, n3553, n3553, n3554, n3554, n3555, n3555, n3556, n3556,
 n3557, n3557, n3558, n3558, n3559, n3559, n3560, n3560, n3561, n3561, n3562, n3562, n3563, n3563, n3564, n3564, n3565, n3565, n3566, n3566,
 n3567, n3567, n3568, n3568, n3569, n3569, n3570, n3570, n3571, n3571, n3572, n3572, n3573, n3573, n3574, n3574, n3575, n3575, n3576, n3576,
 n3577, n3577, n3578, n3578, n3579, n3579, n3580, n3580, n3581, n3581, n3582, n3582, n3583, n3583, n3584, n3584, n3585, n3585, n3586, n3586,
 n3587, n3587, n3588;

 OR2X1TS U1658 ( .A(n3556), .A(n3556_n), .B(n3563), .B(n3563_n), .Y(n3202_n), .Y(n3202) );
 NOR2X1TS U1659 ( .A(n2716), .A(n2716_n), .B(n2819), .B(n2819_n), .Y(n2617_n), .Y(n2617) );
 NAND2X1TS U1660 ( .A(n2851), .A(n2851_n), .B(n2744), .B(n2744_n), .Y(n2618_n), .Y(n2618) );
 NAND2X1TS U1661 ( .A(n3391), .A(n3391_n), .B(n2618), .B(n2618_n), .Y(n2619_n), .Y(n2619) );
 NOR2X1TS U1662 ( .A(n2617), .A(n2617_n), .B(n2619), .B(n2619_n), .Y(n2620_n), .Y(n2620) );
 NAND2X1TS U1663 ( .A(n3018), .A(n3018_n), .B(n2620), .B(n2620_n), .Y(n2621_n), .Y(n2621) );
 NOR2X1TS U1664 ( .A(n2838), .A(n2838_n), .B(n2774), .B(n2774_n), .Y(n2622_n), .Y(n2622) );
 NOR2X1TS U1665 ( .A(n2771), .A(n2771_n), .B(n2768), .B(n2768_n), .Y(n2623_n), .Y(n2623) );
 NOR2X1TS U1666 ( .A(n3222), .A(n3222_n), .B(n2704), .B(n2704_n), .Y(n2624_n), .Y(n2624) );
 NOR2X1TS U1667 ( .A(n2782), .A(n2782_n), .B(n2815), .B(n2815_n), .Y(n2625_n), .Y(n2625) );
 NOR2X1TS U1668 ( .A(n2622), .A(n2622_n), .B(n2623), .B(n2623_n), .Y(n2626_n), .Y(n2626) );
 NOR2X1TS U1669 ( .A(n2624), .A(n2624_n), .B(n2625), .B(n2625_n), .Y(n2627_n), .Y(n2627) );
 NAND2X1TS U1670 ( .A(n2626), .A(n2626_n), .B(n2627), .B(n2627_n), .Y(n2628_n), .Y(n2628) );
 NOR2X1TS U1671 ( .A(n3357), .A(n3357_n), .B(n3358), .B(n3358_n), .Y(n2629_n), .Y(n2629) );
 NAND2X1TS U1672 ( .A(n3085), .A(n3085_n), .B(n3356), .B(n3356_n), .Y(n2630_n), .Y(n2630) );
 NAND2X1TS U1673 ( .A(n2629), .A(n2629_n), .B(n2630), .B(n2630_n), .Y(n2631_n), .Y(n2631) );
 NOR2X1TS U1674 ( .A(n2628), .A(n2628_n), .B(n2631), .B(n2631_n), .Y(n2632_n), .Y(n2632) );
 NAND2X1TS U1675 ( .A(n3017), .A(n3017_n), .B(n2632), .B(n2632_n), .Y(n2633_n), .Y(n2633) );
 NOR2X1TS U1676 ( .A(n2621), .A(n2621_n), .B(n2633), .B(n2633_n), .Y(n2634_n), .Y(n2634) );
 NAND2X1TS U1677 ( .A(n2965), .A(n2965_n), .B(n2634), .B(n2634_n), .Y(n2635_n), .Y(n2635) );
 NOR2BX1TS U1678 ( .AN(n2955), .AN(n2955_n), .B(n2635), .B(n2635_n), .Y(n3060_n), .Y(n3060) );
 NAND2X1TS U1679 ( .A(n2877), .A(n2877_n), .B(n2784), .B(n2784_n), .Y(n2636_n), .Y(n2636) );
 NAND2X1TS U1680 ( .A(n3391), .A(n3391_n), .B(n2636), .B(n2636_n), .Y(n2637_n), .Y(n2637) );
 NOR2X1TS U1681 ( .A(n3462), .A(n3462_n), .B(n3463), .B(n3463_n), .Y(n2638_n), .Y(n2638) );
 NOR2X1TS U1682 ( .A(n2894), .A(n2894_n), .B(n3461), .B(n3461_n), .Y(n2639_n), .Y(n2639) );
 NAND2X1TS U1683 ( .A(n2871), .A(n2871_n), .B(n2639), .B(n2639_n), .Y(n2640_n), .Y(n2640) );
 NAND2X1TS U1684 ( .A(n2638), .A(n2638_n), .B(n2640), .B(n2640_n), .Y(n2641_n), .Y(n2641) );
 NAND2X1TS U1685 ( .A(n3004), .A(n3004_n), .B(n3458), .B(n3458_n), .Y(n2642_n), .Y(n2642) );
 NAND2X1TS U1686 ( .A(n3114), .A(n3114_n), .B(n2642), .B(n2642_n), .Y(n2643_n), .Y(n2643) );
 NOR2X1TS U1687 ( .A(n2831), .A(n2831_n), .B(n2982), .B(n2982_n), .Y(n2644_n), .Y(n2644) );
 NOR2X1TS U1688 ( .A(n2788), .A(n2788_n), .B(n2990), .B(n2990_n), .Y(n2645_n), .Y(n2645) );
 NOR2X1TS U1689 ( .A(n2641), .A(n2641_n), .B(n2643), .B(n2643_n), .Y(n2646_n), .Y(n2646) );
 NOR2X1TS U1690 ( .A(n2644), .A(n2644_n), .B(n2645), .B(n2645_n), .Y(n2647_n), .Y(n2647) );
 NAND2X1TS U1691 ( .A(n2646), .A(n2646_n), .B(n2647), .B(n2647_n), .Y(n2648_n), .Y(n2648) );
 NOR2X1TS U1692 ( .A(n2794), .A(n2794_n), .B(n3095), .B(n3095_n), .Y(n2649_n), .Y(n2649) );
 NOR2X1TS U1693 ( .A(n2637), .A(n2637_n), .B(n2648), .B(n2648_n), .Y(n2650_n), .Y(n2650) );
 NOR2X1TS U1694 ( .A(n3176), .A(n3176_n), .B(n2649), .B(n2649_n), .Y(n2651_n), .Y(n2651) );
 NAND2X1TS U1695 ( .A(n2650), .A(n2650_n), .B(n2651), .B(n2651_n), .Y(n2652_n), .Y(n2652) );
 NAND2BX1TS U1696 ( .AN(n2652), .AN(n2652_n), .B(n3248), .B(n3248_n), .Y(n2653_n), .Y(n2653) );
 NOR2X1TS U1697 ( .A(n3053), .A(n3053_n), .B(n2653), .B(n2653_n), .Y(n2654_n), .Y(n2654) );
 NAND2X1TS U1698 ( .A(n3164), .A(n3164_n), .B(n2654), .B(n2654_n), .Y(d[0]_n), .Y(d[0]) );
 AND2X1TS U1699 ( .A(n3428), .A(n3428_n), .B(n3500), .B(n3500_n), .Y(n3141_n), .Y(n3141) );
 NOR2BX1TS U1700 ( .AN(n3248), .AN(n3248_n), .B(n3165), .B(n3165_n), .Y(n2655_n), .Y(n2655) );
 NAND2X1TS U1701 ( .A(n2787), .A(n2787_n), .B(n2778), .B(n2778_n), .Y(n2656_n), .Y(n2656) );
 NAND2X1TS U1702 ( .A(n3115), .A(n3115_n), .B(n2737), .B(n2737_n), .Y(n2657_n), .Y(n2657) );
 NAND2X1TS U1703 ( .A(n2656), .A(n2656_n), .B(n2657), .B(n2657_n), .Y(n2658_n), .Y(n2658) );
 NAND2X1TS U1704 ( .A(n3220), .A(n3220_n), .B(n3219), .B(n3219_n), .Y(n2659_n), .Y(n2659) );
 NOR2X1TS U1705 ( .A(n3223), .A(n3223_n), .B(n3224), .B(n3224_n), .Y(n2660_n), .Y(n2660) );
 NAND2X1TS U1706 ( .A(n2745), .A(n2745_n), .B(n3221), .B(n3221_n), .Y(n2661_n), .Y(n2661) );
 NAND2X1TS U1707 ( .A(n2660), .A(n2660_n), .B(n2661), .B(n2661_n), .Y(n2662_n), .Y(n2662) );
 NOR2X1TS U1708 ( .A(n2833), .A(n2833_n), .B(n2807), .B(n2807_n), .Y(n2663_n), .Y(n2663) );
 AND2X1TS U1709 ( .A(n2846), .A(n2846_n), .B(n2748), .B(n2748_n), .Y(n2664_n), .Y(n2664) );
 NOR2X1TS U1710 ( .A(n2659), .A(n2659_n), .B(n2662), .B(n2662_n), .Y(n2665_n), .Y(n2665) );
 NOR2X1TS U1711 ( .A(n2663), .A(n2663_n), .B(n2664), .B(n2664_n), .Y(n2666_n), .Y(n2666) );
 NAND2X1TS U1712 ( .A(n2665), .A(n2665_n), .B(n2666), .B(n2666_n), .Y(n2667_n), .Y(n2667) );
 NOR2X1TS U1713 ( .A(n2658), .A(n2658_n), .B(n2667), .B(n2667_n), .Y(n2668_n), .Y(n2668) );
 NAND2X1TS U1714 ( .A(n3031), .A(n3031_n), .B(n2668), .B(n2668_n), .Y(n2669_n), .Y(n2669) );
 NOR2X1TS U1715 ( .A(n2669), .A(n2669_n), .B(n3179), .B(n3179_n), .Y(n2670_n), .Y(n2670) );
 NOR2X1TS U1716 ( .A(n3196), .A(n3196_n), .B(n3203), .B(n3203_n), .Y(n2671_n), .Y(n2671) );
 NAND2X1TS U1717 ( .A(n2670), .A(n2670_n), .B(n2671), .B(n2671_n), .Y(n2672_n), .Y(n2672) );
 NOR2X1TS U1718 ( .A(n3247), .A(n3247_n), .B(n2672), .B(n2672_n), .Y(n2673_n), .Y(n2673) );
 NAND2X1TS U1719 ( .A(n2655), .A(n2655_n), .B(n2673), .B(n2673_n), .Y(d[2]_n), .Y(d[2]) );
 NOR2X1TS U1720 ( .A(n2840), .A(n2840_n), .B(n3171), .B(n3171_n), .Y(n2674_n), .Y(n2674) );
 NOR2X1TS U1721 ( .A(n2830), .A(n2830_n), .B(n2712), .B(n2712_n), .Y(n2675_n), .Y(n2675) );
 NOR2X1TS U1722 ( .A(n2674), .A(n2674_n), .B(n2675), .B(n2675_n), .Y(n2676_n), .Y(n2676) );
 NAND2X1TS U1723 ( .A(n2851), .A(n2851_n), .B(n2779), .B(n2779_n), .Y(n2677_n), .Y(n2677) );
 NAND2X1TS U1724 ( .A(n2676), .A(n2676_n), .B(n2677), .B(n2677_n), .Y(n2678_n), .Y(n2678) );
 NAND2X1TS U1725 ( .A(n2726), .A(n2726_n), .B(n3170), .B(n3170_n), .Y(n2679_n), .Y(n2679) );
 NAND2X1TS U1726 ( .A(n2785), .A(n2785_n), .B(n3166), .B(n3166_n), .Y(n2680_n), .Y(n2680) );
 NAND2X1TS U1727 ( .A(n2679), .A(n2679_n), .B(n2680), .B(n2680_n), .Y(n2681_n), .Y(n2681) );
 NOR2BX1TS U1728 ( .AN(n2849), .AN(n2849_n), .B(n3167), .B(n3167_n), .Y(n2682_n), .Y(n2682) );
 NOR2X1TS U1729 ( .A(n2682), .A(n2682_n), .B(n2681), .B(n2681_n), .Y(n2683_n), .Y(n2683) );
 NAND2X1TS U1730 ( .A(n2933), .A(n2933_n), .B(n3168), .B(n3168_n), .Y(n2684_n), .Y(n2684) );
 NAND2X1TS U1731 ( .A(n2683), .A(n2683_n), .B(n2684), .B(n2684_n), .Y(n2685_n), .Y(n2685) );
 NOR2X1TS U1732 ( .A(n2719), .A(n2719_n), .B(n2761), .B(n2761_n), .Y(n2686_n), .Y(n2686) );
 NOR2X1TS U1733 ( .A(n3172), .A(n3172_n), .B(n2686), .B(n2686_n), .Y(n2687_n), .Y(n2687) );
 NAND2X1TS U1734 ( .A(n3070), .A(n3070_n), .B(n2687), .B(n2687_n), .Y(n2688_n), .Y(n2688) );
 NOR2X1TS U1735 ( .A(n2678), .A(n2678_n), .B(n2685), .B(n2685_n), .Y(n2689_n), .Y(n2689) );
 NOR2X1TS U1736 ( .A(n2688), .A(n2688_n), .B(n3165), .B(n3165_n), .Y(n2690_n), .Y(n2690) );
 NAND2X1TS U1737 ( .A(n2689), .A(n2689_n), .B(n2690), .B(n2690_n), .Y(n2691_n), .Y(n2691) );
 NOR2X1TS U1738 ( .A(n3028), .A(n3028_n), .B(n2691), .B(n2691_n), .Y(n2692_n), .Y(n2692) );
 NAND2X1TS U1739 ( .A(n3164), .A(n3164_n), .B(n2692), .B(n2692_n), .Y(d[3]_n), .Y(d[3]) );
 AND2X2TS U1740 ( .A(n3500), .A(n3500_n), .B(n3555), .B(n3555_n), .Y(n2693_n), .Y(n2693) );
 AND2X2TS U1741 ( .A(n2706), .A(n2706_n), .B(n3555), .B(n3555_n), .Y(n2694_n), .Y(n2694) );
 AND2X2TS U1742 ( .A(n3500), .A(n3500_n), .B(n3460), .B(n3460_n), .Y(n2695_n), .Y(n2695) );
 AND2X2TS U1743 ( .A(n2913), .A(n2913_n), .B(n3446), .B(n3446_n), .Y(n2696_n), .Y(n2696) );
 OR2X2TS U1744 ( .A(n3568), .A(n3568_n), .B(n3569), .B(n3569_n), .Y(n2697_n), .Y(n2697) );
 AND2X2TS U1745 ( .A(n3446), .A(n3446_n), .B(n3562), .B(n3562_n), .Y(n2698_n), .Y(n2698) );
 AND2X2TS U1746 ( .A(n2903), .A(n2903_n), .B(n3304), .B(n3304_n), .Y(n2699_n), .Y(n2699) );
 AND2X2TS U1747 ( .A(n3499), .A(n3499_n), .B(n3459), .B(n3459_n), .Y(n2700_n), .Y(n2700) );
 AND2X2TS U1748 ( .A(n3370), .A(n3370_n), .B(n3466), .B(n3466_n), .Y(n2701_n), .Y(n2701) );
 OR2X2TS U1749 ( .A(n2863), .A(n2863_n), .B(n2857), .B(n2857_n), .Y(n2702_n), .Y(n2702) );
 NAND2X1TS U1750 ( .A(n2905), .A(n2905_n), .B(n2893), .B(n2893_n), .Y(n2703_n), .Y(n2703) );
 INVXLTS U1751 ( .A(n2994), .A(n2994_n), .Y(n2704_n), .Y(n2704) );
 INVXLTS U1752 ( .A(n2994), .A(n2994_n), .Y(n2705_n), .Y(n2705) );
 INVXLTS U1753 ( .A(n2703), .A(n2703_n), .Y(n2706_n), .Y(n2706) );
 INVXLTS U1754 ( .A(n2703), .A(n2703_n), .Y(n2707_n), .Y(n2707) );
 INVXLTS U1755 ( .A(n3460), .A(n3460_n), .Y(n2708_n), .Y(n2708) );
 INVXLTS U1756 ( .A(n2708), .A(n2708_n), .Y(n2709_n), .Y(n2709) );
 INVXLTS U1757 ( .A(n2933), .A(n2933_n), .Y(n2710_n), .Y(n2710) );
 INVXLTS U1758 ( .A(n2702), .A(n2702_n), .Y(n2711_n), .Y(n2711) );
 INVXLTS U1759 ( .A(n2702), .A(n2702_n), .Y(n2712_n), .Y(n2712) );
 INVXLTS U1760 ( .A(n3096), .A(n3096_n), .Y(n2713_n), .Y(n2713) );
 INVXLTS U1761 ( .A(n3096), .A(n3096_n), .Y(n2714_n), .Y(n2714) );
 INVXLTS U1762 ( .A(n2939), .A(n2939_n), .Y(n2715_n), .Y(n2715) );
 INVXLTS U1763 ( .A(n2939), .A(n2939_n), .Y(n2716_n), .Y(n2716) );
 INVXLTS U1764 ( .A(n3131), .A(n3131_n), .Y(n2717_n), .Y(n2717) );
 INVXLTS U1765 ( .A(n3131), .A(n3131_n), .Y(n2718_n), .Y(n2718) );
 INVXLTS U1766 ( .A(n2925), .A(n2925_n), .Y(n2719_n), .Y(n2719) );
 INVXLTS U1767 ( .A(n2925), .A(n2925_n), .Y(n2720_n), .Y(n2720) );
 INVXLTS U1768 ( .A(n2975), .A(n2975_n), .Y(n2721_n), .Y(n2721) );
 INVXLTS U1769 ( .A(n2975), .A(n2975_n), .Y(n2722_n), .Y(n2722) );
 INVXLTS U1770 ( .A(n2700), .A(n2700_n), .Y(n2723_n), .Y(n2723) );
 INVXLTS U1771 ( .A(n2700), .A(n2700_n), .Y(n2724_n), .Y(n2724) );
 INVXLTS U1772 ( .A(n3202), .A(n3202_n), .Y(n2725_n), .Y(n2725) );
 INVXLTS U1773 ( .A(n3202), .A(n3202_n), .Y(n2726_n), .Y(n2726) );
 INVXLTS U1774 ( .A(n2935), .A(n2935_n), .Y(n2727_n), .Y(n2727) );
 INVXLTS U1775 ( .A(n2935), .A(n2935_n), .Y(n2728_n), .Y(n2728) );
 INVXLTS U1776 ( .A(n2697), .A(n2697_n), .Y(n2729_n), .Y(n2729) );
 INVXLTS U1777 ( .A(n2697), .A(n2697_n), .Y(n2730_n), .Y(n2730) );
 INVXLTS U1778 ( .A(n2699), .A(n2699_n), .Y(n2731_n), .Y(n2731) );
 INVXLTS U1779 ( .A(n2699), .A(n2699_n), .Y(n2732_n), .Y(n2732) );
 INVXLTS U1780 ( .A(n2698), .A(n2698_n), .Y(n2733_n), .Y(n2733) );
 INVXLTS U1781 ( .A(n2698), .A(n2698_n), .Y(n2734_n), .Y(n2734) );
 INVXLTS U1782 ( .A(n3161), .A(n3161_n), .Y(n2735_n), .Y(n2735) );
 INVXLTS U1783 ( .A(n3161), .A(n3161_n), .Y(n2736_n), .Y(n2736) );
 INVXLTS U1784 ( .A(n3080), .A(n3080_n), .Y(n2737_n), .Y(n2737) );
 INVXLTS U1785 ( .A(n3080), .A(n3080_n), .Y(n2738_n), .Y(n2738) );
 INVXLTS U1786 ( .A(n2701), .A(n2701_n), .Y(n2739_n), .Y(n2739) );
 INVXLTS U1787 ( .A(n2701), .A(n2701_n), .Y(n2740_n), .Y(n2740) );
 INVXLTS U1788 ( .A(n2945), .A(n2945_n), .Y(n2741_n), .Y(n2741) );
 INVXLTS U1789 ( .A(n2741), .A(n2741_n), .Y(n2742_n), .Y(n2742) );
 INVXLTS U1790 ( .A(n2741), .A(n2741_n), .Y(n2743_n), .Y(n2743) );
 INVXLTS U1791 ( .A(n2945), .A(n2945_n), .Y(n2744_n), .Y(n2744) );
 INVXLTS U1792 ( .A(n2945), .A(n2945_n), .Y(n2745_n), .Y(n2745) );
 INVXLTS U1793 ( .A(n3006), .A(n3006_n), .Y(n2746_n), .Y(n2746) );
 INVXLTS U1794 ( .A(n2746), .A(n2746_n), .Y(n2747_n), .Y(n2747) );
 INVXLTS U1795 ( .A(n2746), .A(n2746_n), .Y(n2748_n), .Y(n2748) );
 INVXLTS U1796 ( .A(n3023), .A(n3023_n), .Y(n2749_n), .Y(n2749) );
 INVXLTS U1797 ( .A(n2749), .A(n2749_n), .Y(n2750_n), .Y(n2750) );
 INVXLTS U1798 ( .A(n2988), .A(n2988_n), .Y(n2751_n), .Y(n2751) );
 INVXLTS U1799 ( .A(n2751), .A(n2751_n), .Y(n2752_n), .Y(n2752) );
 INVXLTS U1800 ( .A(n2751), .A(n2751_n), .Y(n2753_n), .Y(n2753) );
 INVXLTS U1801 ( .A(n3089), .A(n3089_n), .Y(n2754_n), .Y(n2754) );
 INVXLTS U1802 ( .A(n3089), .A(n3089_n), .Y(n2756_n), .Y(n2756) );
 INVXLTS U1803 ( .A(n3089), .A(n3089_n), .Y(n2755_n), .Y(n2755) );
 INVXLTS U1804 ( .A(n2928), .A(n2928_n), .Y(n2757_n), .Y(n2757) );
 INVXLTS U1805 ( .A(n2928), .A(n2928_n), .Y(n2759_n), .Y(n2759) );
 INVXLTS U1806 ( .A(n2928), .A(n2928_n), .Y(n2758_n), .Y(n2758) );
 INVXLTS U1807 ( .A(n2693), .A(n2693_n), .Y(n2760_n), .Y(n2760) );
 INVXLTS U1808 ( .A(n2693), .A(n2693_n), .Y(n2762_n), .Y(n2762) );
 INVXLTS U1809 ( .A(n2693), .A(n2693_n), .Y(n2761_n), .Y(n2761) );
 INVXLTS U1810 ( .A(n3125), .A(n3125_n), .Y(n2763_n), .Y(n2763) );
 INVXLTS U1811 ( .A(n3125), .A(n3125_n), .Y(n2765_n), .Y(n2765) );
 INVXLTS U1812 ( .A(n3125), .A(n3125_n), .Y(n2764_n), .Y(n2764) );
 INVXLTS U1813 ( .A(n2986), .A(n2986_n), .Y(n2766_n), .Y(n2766) );
 INVXLTS U1814 ( .A(n2986), .A(n2986_n), .Y(n2768_n), .Y(n2768) );
 INVXLTS U1815 ( .A(n2986), .A(n2986_n), .Y(n2767_n), .Y(n2767) );
 INVXLTS U1816 ( .A(n2760), .A(n2760_n), .Y(n2769_n), .Y(n2769) );
 INVXLTS U1817 ( .A(n2762), .A(n2762_n), .Y(n2770_n), .Y(n2770) );
 INVXLTS U1818 ( .A(n3051), .A(n3051_n), .Y(n2772_n), .Y(n2772) );
 INVXLTS U1819 ( .A(n3051), .A(n3051_n), .Y(n2771_n), .Y(n2771) );
 INVXLTS U1820 ( .A(n3013), .A(n3013_n), .Y(n2773_n), .Y(n2773) );
 INVXLTS U1821 ( .A(n2773), .A(n2773_n), .Y(n2774_n), .Y(n2774) );
 INVXLTS U1822 ( .A(n2773), .A(n2773_n), .Y(n2776_n), .Y(n2776) );
 INVXLTS U1823 ( .A(n2773), .A(n2773_n), .Y(n2775_n), .Y(n2775) );
 INVXLTS U1824 ( .A(n3085), .A(n3085_n), .Y(n2777_n), .Y(n2777) );
 INVXLTS U1825 ( .A(n2777), .A(n2777_n), .Y(n2778_n), .Y(n2778) );
 INVXLTS U1826 ( .A(n2777), .A(n2777_n), .Y(n2779_n), .Y(n2779) );
 INVXLTS U1827 ( .A(n3077), .A(n3077_n), .Y(n2780_n), .Y(n2780) );
 INVXLTS U1828 ( .A(n3077), .A(n3077_n), .Y(n2782_n), .Y(n2782) );
 INVXLTS U1829 ( .A(n3077), .A(n3077_n), .Y(n2781_n), .Y(n2781) );
 INVXLTS U1830 ( .A(n2791), .A(n2791_n), .Y(n2783_n), .Y(n2783) );
 INVXLTS U1831 ( .A(n2793), .A(n2793_n), .Y(n2784_n), .Y(n2784) );
 INVXLTS U1832 ( .A(n3013), .A(n3013_n), .Y(n2785_n), .Y(n2785) );
 INVXLTS U1833 ( .A(n3013), .A(n3013_n), .Y(n2787_n), .Y(n2787) );
 INVXLTS U1834 ( .A(n3013), .A(n3013_n), .Y(n2786_n), .Y(n2786) );
 INVXLTS U1835 ( .A(n2763), .A(n2763_n), .Y(n2788_n), .Y(n2788) );
 INVXLTS U1836 ( .A(n2765), .A(n2765_n), .Y(n2790_n), .Y(n2790) );
 INVXLTS U1837 ( .A(n2764), .A(n2764_n), .Y(n2789_n), .Y(n2789) );
 INVXLTS U1838 ( .A(n2695), .A(n2695_n), .Y(n2791_n), .Y(n2791) );
 INVXLTS U1839 ( .A(n2695), .A(n2695_n), .Y(n2793_n), .Y(n2793) );
 INVXLTS U1840 ( .A(n2695), .A(n2695_n), .Y(n2792_n), .Y(n2792) );
 INVXLTS U1841 ( .A(n2694), .A(n2694_n), .Y(n2794_n), .Y(n2794) );
 INVXLTS U1842 ( .A(n2694), .A(n2694_n), .Y(n2796_n), .Y(n2796) );
 INVXLTS U1843 ( .A(n2694), .A(n2694_n), .Y(n2795_n), .Y(n2795) );
 INVXLTS U1844 ( .A(n2988), .A(n2988_n), .Y(n2798_n), .Y(n2798) );
 INVXLTS U1845 ( .A(n2988), .A(n2988_n), .Y(n2797_n), .Y(n2797) );
 INVXLTS U1846 ( .A(n3015), .A(n3015_n), .Y(n2799_n), .Y(n2799) );
 INVXLTS U1847 ( .A(n2799), .A(n2799_n), .Y(n2800_n), .Y(n2800) );
 INVXLTS U1848 ( .A(n2799), .A(n2799_n), .Y(n2801_n), .Y(n2801) );
 INVXLTS U1849 ( .A(n3141), .A(n3141_n), .Y(n2802_n), .Y(n2802) );
 INVXLTS U1850 ( .A(n3141), .A(n3141_n), .Y(n2804_n), .Y(n2804) );
 INVXLTS U1851 ( .A(n3141), .A(n3141_n), .Y(n2803_n), .Y(n2803) );
 INVXLTS U1852 ( .A(n2946), .A(n2946_n), .Y(n2805_n), .Y(n2805) );
 INVXLTS U1853 ( .A(n2946), .A(n2946_n), .Y(n2807_n), .Y(n2807) );
 INVXLTS U1854 ( .A(n2946), .A(n2946_n), .Y(n2806_n), .Y(n2806) );
 INVXLTS U1855 ( .A(n2699), .A(n2699_n), .Y(n2808_n), .Y(n2808) );
 INVXLTS U1856 ( .A(n2808), .A(n2808_n), .Y(n2809_n), .Y(n2809) );
 INVXLTS U1857 ( .A(n2808), .A(n2808_n), .Y(n2811_n), .Y(n2811) );
 INVXLTS U1858 ( .A(n2808), .A(n2808_n), .Y(n2810_n), .Y(n2810) );
 INVXLTS U1859 ( .A(n3096), .A(n3096_n), .Y(n2812_n), .Y(n2812) );
 INVXLTS U1860 ( .A(n2812), .A(n2812_n), .Y(n2813_n), .Y(n2813) );
 INVXLTS U1861 ( .A(n2812), .A(n2812_n), .Y(n2815_n), .Y(n2815) );
 INVXLTS U1862 ( .A(n2812), .A(n2812_n), .Y(n2814_n), .Y(n2814) );
 INVXLTS U1863 ( .A(n2796), .A(n2796_n), .Y(n2816_n), .Y(n2816) );
 INVXLTS U1864 ( .A(n2794), .A(n2794_n), .Y(n2817_n), .Y(n2817) );
 INVXLTS U1865 ( .A(n3131), .A(n3131_n), .Y(n2818_n), .Y(n2818) );
 INVXLTS U1866 ( .A(n2818), .A(n2818_n), .Y(n2819_n), .Y(n2819) );
 INVXLTS U1867 ( .A(n2818), .A(n2818_n), .Y(n2821_n), .Y(n2821) );
 INVXLTS U1868 ( .A(n2818), .A(n2818_n), .Y(n2820_n), .Y(n2820) );
 INVXLTS U1869 ( .A(n2696), .A(n2696_n), .Y(n2822_n), .Y(n2822) );
 INVXLTS U1870 ( .A(n2696), .A(n2696_n), .Y(n2824_n), .Y(n2824) );
 INVXLTS U1871 ( .A(n2696), .A(n2696_n), .Y(n2823_n), .Y(n2823) );
 INVXLTS U1872 ( .A(n3080), .A(n3080_n), .Y(n2825_n), .Y(n2825) );
 INVXLTS U1873 ( .A(n2825), .A(n2825_n), .Y(n2826_n), .Y(n2826) );
 INVXLTS U1874 ( .A(n2825), .A(n2825_n), .Y(n2828_n), .Y(n2828) );
 INVXLTS U1875 ( .A(n2825), .A(n2825_n), .Y(n2827_n), .Y(n2827) );
 INVXLTS U1876 ( .A(n2755), .A(n2755_n), .Y(n2829_n), .Y(n2829) );
 INVXLTS U1877 ( .A(n2756), .A(n2756_n), .Y(n2830_n), .Y(n2830) );
 INVXLTS U1878 ( .A(n2754), .A(n2754_n), .Y(n2831_n), .Y(n2831) );
 INVXLTS U1879 ( .A(n3202), .A(n3202_n), .Y(n2832_n), .Y(n2832) );
 INVXLTS U1880 ( .A(n2832), .A(n2832_n), .Y(n2835_n), .Y(n2835) );
 INVXLTS U1881 ( .A(n2832), .A(n2832_n), .Y(n2833_n), .Y(n2833) );
 INVXLTS U1882 ( .A(n2832), .A(n2832_n), .Y(n2834_n), .Y(n2834) );
 INVXLTS U1883 ( .A(n2954), .A(n2954_n), .Y(n2836_n), .Y(n2836) );
 INVXLTS U1884 ( .A(n2836), .A(n2836_n), .Y(n2837_n), .Y(n2837) );
 INVXLTS U1885 ( .A(n2836), .A(n2836_n), .Y(n2838_n), .Y(n2838) );
 INVXLTS U1886 ( .A(n2836), .A(n2836_n), .Y(n2839_n), .Y(n2839) );
 INVXLTS U1887 ( .A(n3051), .A(n3051_n), .Y(n2840_n), .Y(n2840) );
 INVXLTS U1888 ( .A(n2840), .A(n2840_n), .Y(n2841_n), .Y(n2841) );
 INVXLTS U1889 ( .A(n2840), .A(n2840_n), .Y(n2842_n), .Y(n2842) );
 INVXLTS U1890 ( .A(n2700), .A(n2700_n), .Y(n2843_n), .Y(n2843) );
 INVXLTS U1891 ( .A(n2843), .A(n2843_n), .Y(n2844_n), .Y(n2844) );
 INVXLTS U1892 ( .A(n2843), .A(n2843_n), .Y(n2846_n), .Y(n2846) );
 INVXLTS U1893 ( .A(n2843), .A(n2843_n), .Y(n2845_n), .Y(n2845) );
 INVXLTS U1894 ( .A(n2946), .A(n2946_n), .Y(n2847_n), .Y(n2847) );
 INVXLTS U1895 ( .A(n2847), .A(n2847_n), .Y(n2848_n), .Y(n2848) );
 INVXLTS U1896 ( .A(n2847), .A(n2847_n), .Y(n2849_n), .Y(n2849) );
 INVXLTS U1897 ( .A(n3141), .A(n3141_n), .Y(n2850_n), .Y(n2850) );
 INVXLTS U1898 ( .A(n2850), .A(n2850_n), .Y(n2851_n), .Y(n2851) );
 INVXLTS U1899 ( .A(n2850), .A(n2850_n), .Y(n2852_n), .Y(n2852) );
 INVXLTS U1900 ( .A(n3161), .A(n3161_n), .Y(n2853_n), .Y(n2853) );
 INVXLTS U1901 ( .A(n2853), .A(n2853_n), .Y(n2854_n), .Y(n2854) );
 INVXLTS U1902 ( .A(n2853), .A(n2853_n), .Y(n2855_n), .Y(n2855) );
 INVXLTS U1903 ( .A(n2939), .A(n2939_n), .Y(n2856_n), .Y(n2856) );
 INVXLTS U1904 ( .A(n2856), .A(n2856_n), .Y(n2857_n), .Y(n2857) );
 INVXLTS U1905 ( .A(n2856), .A(n2856_n), .Y(n2858_n), .Y(n2858) );
 INVXLTS U1906 ( .A(n2767), .A(n2767_n), .Y(n2859_n), .Y(n2859) );
 INVXLTS U1907 ( .A(n2766), .A(n2766_n), .Y(n2860_n), .Y(n2860) );
 INVXLTS U1908 ( .A(n2933), .A(n2933_n), .Y(n2861_n), .Y(n2861) );
 INVXLTS U1909 ( .A(n2861), .A(n2861_n), .Y(n2862_n), .Y(n2862) );
 INVXLTS U1910 ( .A(n2861), .A(n2861_n), .Y(n2863_n), .Y(n2863) );
 INVXLTS U1911 ( .A(n3077), .A(n3077_n), .Y(n2864_n), .Y(n2864) );
 INVXLTS U1912 ( .A(n2864), .A(n2864_n), .Y(n2865_n), .Y(n2865) );
 INVXLTS U1913 ( .A(n2864), .A(n2864_n), .Y(n2867_n), .Y(n2867) );
 INVXLTS U1914 ( .A(n2864), .A(n2864_n), .Y(n2866_n), .Y(n2866) );
 INVXLTS U1915 ( .A(n2975), .A(n2975_n), .Y(n2868_n), .Y(n2868) );
 INVXLTS U1916 ( .A(n2868), .A(n2868_n), .Y(n2869_n), .Y(n2869) );
 INVXLTS U1917 ( .A(n2868), .A(n2868_n), .Y(n2871_n), .Y(n2871) );
 INVXLTS U1918 ( .A(n2868), .A(n2868_n), .Y(n2870_n), .Y(n2870) );
 INVXLTS U1919 ( .A(n2994), .A(n2994_n), .Y(n2872_n), .Y(n2872) );
 INVXLTS U1920 ( .A(n2872), .A(n2872_n), .Y(n2873_n), .Y(n2873) );
 INVXLTS U1921 ( .A(n2872), .A(n2872_n), .Y(n2874_n), .Y(n2874) );
 INVXLTS U1922 ( .A(n2872), .A(n2872_n), .Y(n2875_n), .Y(n2875) );
 INVXLTS U1923 ( .A(n2928), .A(n2928_n), .Y(n2876_n), .Y(n2876) );
 INVXLTS U1924 ( .A(n2876), .A(n2876_n), .Y(n2877_n), .Y(n2877) );
 INVXLTS U1925 ( .A(n2876), .A(n2876_n), .Y(n2878_n), .Y(n2878) );
 INVXLTS U1926 ( .A(n2876), .A(n2876_n), .Y(n2879_n), .Y(n2879) );
 INVXLTS U1927 ( .A(n2925), .A(n2925_n), .Y(n2880_n), .Y(n2880) );
 INVXLTS U1928 ( .A(n2880), .A(n2880_n), .Y(n2881_n), .Y(n2881) );
 INVXLTS U1929 ( .A(n2880), .A(n2880_n), .Y(n2882_n), .Y(n2882) );
 INVXLTS U1930 ( .A(n2880), .A(n2880_n), .Y(n2883_n), .Y(n2883) );
 INVXLTS U1931 ( .A(n2935), .A(n2935_n), .Y(n2884_n), .Y(n2884) );
 INVXLTS U1932 ( .A(n2884), .A(n2884_n), .Y(n2885_n), .Y(n2885) );
 INVXLTS U1933 ( .A(n2884), .A(n2884_n), .Y(n2888_n), .Y(n2888) );
 INVXLTS U1934 ( .A(n2884), .A(n2884_n), .Y(n2886_n), .Y(n2886) );
 INVXLTS U1935 ( .A(n2884), .A(n2884_n), .Y(n2887_n), .Y(n2887) );
 INVXLTS U1936 ( .A(a[2]), .A(a[2]_n), .Y(n2889_n), .Y(n2889) );
 INVXLTS U1937 ( .A(n2889), .A(n2889_n), .Y(n2890_n), .Y(n2890) );
 INVXLTS U1938 ( .A(n2889), .A(n2889_n), .Y(n2891_n), .Y(n2891) );
 INVXLTS U1939 ( .A(a[7]), .A(a[7]_n), .Y(n2892_n), .Y(n2892) );
 INVXLTS U1940 ( .A(n2892), .A(n2892_n), .Y(n2893_n), .Y(n2893) );
 INVXLTS U1941 ( .A(n2892), .A(n2892_n), .Y(n2894_n), .Y(n2894) );
 INVXLTS U1942 ( .A(a[6]), .A(a[6]_n), .Y(n2895_n), .Y(n2895) );
 INVXLTS U1943 ( .A(n2895), .A(n2895_n), .Y(n2896_n), .Y(n2896) );
 INVXLTS U1944 ( .A(n2895), .A(n2895_n), .Y(n2897_n), .Y(n2897) );
 INVXLTS U1945 ( .A(a[3]), .A(a[3]_n), .Y(n2898_n), .Y(n2898) );
 INVXLTS U1946 ( .A(n2898), .A(n2898_n), .Y(n2899_n), .Y(n2899) );
 INVXLTS U1947 ( .A(n2898), .A(n2898_n), .Y(n2900_n), .Y(n2900) );
 INVXLTS U1948 ( .A(a[0]), .A(a[0]_n), .Y(n2901_n), .Y(n2901) );
 INVXLTS U1949 ( .A(n2901), .A(n2901_n), .Y(n2902_n), .Y(n2902) );
 INVXLTS U1950 ( .A(n2901), .A(n2901_n), .Y(n2903_n), .Y(n2903) );
 INVXLTS U1951 ( .A(a[5]), .A(a[5]_n), .Y(n2904_n), .Y(n2904) );
 INVXLTS U1952 ( .A(n2904), .A(n2904_n), .Y(n2905_n), .Y(n2905) );
 INVXLTS U1953 ( .A(n2904), .A(n2904_n), .Y(n2906_n), .Y(n2906) );
 INVXLTS U1954 ( .A(a[4]), .A(a[4]_n), .Y(n2907_n), .Y(n2907) );
 INVXLTS U1955 ( .A(n2907), .A(n2907_n), .Y(n2908_n), .Y(n2908) );
 INVXLTS U1956 ( .A(n2907), .A(n2907_n), .Y(n2909_n), .Y(n2909) );
 INVXLTS U1957 ( .A(a[1]), .A(a[1]_n), .Y(n2910_n), .Y(n2910) );
 INVXLTS U1958 ( .A(n2910), .A(n2910_n), .Y(n2911_n), .Y(n2911) );
 INVXLTS U1959 ( .A(n2910), .A(n2910_n), .Y(n2913_n), .Y(n2913) );
 INVXLTS U1960 ( .A(n2910), .A(n2910_n), .Y(n2912_n), .Y(n2912) );
 AND2XLTS U1961 ( .A(n2718), .A(n2718_n), .B(n3464), .B(n3464_n), .Y(n3463_n), .Y(n3463) );
 NOR2XLTS U1962 ( .A(n2736), .A(n2736_n), .B(n3465), .B(n3465_n), .Y(n3462_n), .Y(n3462) );
 NOR2XLTS U1963 ( .A(n2963), .A(n2963_n), .B(n2964), .B(n2964_n), .Y(n2962_n), .Y(n2962) );
 NOR2XLTS U1964 ( .A(n2967), .A(n2967_n), .B(n2968), .B(n2968_n), .Y(n2966_n), .Y(n2966) );
 NOR2XLTS U1965 ( .A(n2971), .A(n2971_n), .B(n2972), .B(n2972_n), .Y(n2970_n), .Y(n2970) );
 NOR2XLTS U1966 ( .A(n2977), .A(n2977_n), .B(n2734), .B(n2734_n), .Y(n2971_n), .Y(n2971) );
 NOR2XLTS U1967 ( .A(n2978), .A(n2978_n), .B(n2979), .B(n2979_n), .Y(n2969_n), .Y(n2969) );
 NOR2XLTS U1968 ( .A(n2750), .A(n2750_n), .B(n2745), .B(n2745_n), .Y(n2990_n), .Y(n2990) );
 NOR2XLTS U1969 ( .A(n2917), .A(n2917_n), .B(n2991), .B(n2991_n), .Y(n2961_n), .Y(n2961) );
 NOR2XLTS U1970 ( .A(n3028), .A(n3028_n), .B(n3029), .B(n3029_n), .Y(n3027_n), .Y(n3027) );
 NOR2XLTS U1971 ( .A(n3032), .A(n3032_n), .B(n3033), .B(n3033_n), .Y(n3030_n), .Y(n3030) );
 NOR2XLTS U1972 ( .A(n3036), .A(n3036_n), .B(n3037), .B(n3037_n), .Y(n3035_n), .Y(n3035) );
 NOR2XLTS U1973 ( .A(n2734), .A(n2734_n), .B(n2772), .B(n2772_n), .Y(n3037_n), .Y(n3037) );
 NOR2XLTS U1974 ( .A(n3038), .A(n3038_n), .B(n3039), .B(n3039_n), .Y(n3034_n), .Y(n3034) );
 NOR2XLTS U1975 ( .A(n2711), .A(n2711_n), .B(n2735), .B(n2735_n), .Y(n3039_n), .Y(n3039) );
 NOR2XLTS U1976 ( .A(n3040), .A(n3040_n), .B(n2805), .B(n2805_n), .Y(n3038_n), .Y(n3038) );
 NOR2XLTS U1977 ( .A(n3043), .A(n3043_n), .B(n3044), .B(n3044_n), .Y(n3042_n), .Y(n3042) );
 AND2XLTS U1978 ( .A(n2846), .A(n2846_n), .B(n2976), .B(n2976_n), .Y(n3044_n), .Y(n3044) );
 NOR2XLTS U1979 ( .A(n2891), .A(n2891_n), .B(n2913), .B(n2913_n), .Y(n3046_n), .Y(n3046) );
 NOR2XLTS U1980 ( .A(n3047), .A(n3047_n), .B(n2710), .B(n2710_n), .Y(n3043_n), .Y(n3043) );
 NOR2XLTS U1981 ( .A(n3048), .A(n3048_n), .B(n3049), .B(n3049_n), .Y(n3041_n), .Y(n3041) );
 NOR2XLTS U1982 ( .A(n3050), .A(n3050_n), .B(n2739), .B(n2739_n), .Y(n3049_n), .Y(n3049) );
 NOR2XLTS U1983 ( .A(n2694), .A(n2694_n), .B(n2841), .B(n2841_n), .Y(n3050_n), .Y(n3050) );
 NOR2XLTS U1984 ( .A(n2839), .A(n2839_n), .B(n2947), .B(n2947_n), .Y(n3048_n), .Y(n3048) );
 NOR2XLTS U1985 ( .A(n3052), .A(n3052_n), .B(n3053), .B(n3053_n), .Y(n3026_n), .Y(n3026) );
 OR2XLTS U1986 ( .A(n3203), .A(n3203_n), .B(n3467), .B(n3467_n), .Y(n3053_n), .Y(n3053) );
 NOR2XLTS U1987 ( .A(n3470), .A(n3470_n), .B(n3471), .B(n3471_n), .Y(n3469_n), .Y(n3469) );
 NOR2XLTS U1988 ( .A(n2831), .A(n2831_n), .B(n2824), .B(n2824_n), .Y(n3470_n), .Y(n3470) );
 NOR2XLTS U1989 ( .A(n3474), .A(n3474_n), .B(n3475), .B(n3475_n), .Y(n3468_n), .Y(n3468) );
 NOR2XLTS U1990 ( .A(n3483), .A(n3483_n), .B(n3484), .B(n3484_n), .Y(n3479_n), .Y(n3479) );
 NOR2XLTS U1991 ( .A(n3485), .A(n3485_n), .B(n2821), .B(n2821_n), .Y(n3484_n), .Y(n3484) );
 NOR2XLTS U1992 ( .A(n2858), .A(n2858_n), .B(n2878), .B(n2878_n), .Y(n3485_n), .Y(n3485) );
 NOR2XLTS U1993 ( .A(n3486), .A(n3486_n), .B(n2760), .B(n2760_n), .Y(n3483_n), .Y(n3483) );
 NOR2XLTS U1994 ( .A(n2867), .A(n2867_n), .B(n3446), .B(n3446_n), .Y(n3486_n), .Y(n3486) );
 NOR2XLTS U1995 ( .A(n3056), .A(n3056_n), .B(n3057), .B(n3057_n), .Y(n3055_n), .Y(n3055) );
 NOR2XLTS U1996 ( .A(n2804), .A(n2804_n), .B(n2758), .B(n2758_n), .Y(n3056_n), .Y(n3056) );
 NOR2XLTS U1997 ( .A(n3058), .A(n3058_n), .B(n3059), .B(n3059_n), .Y(n3054_n), .Y(n3054) );
 NOR2XLTS U1998 ( .A(n2963), .A(n2963_n), .B(n3062), .B(n3062_n), .Y(n3061_n), .Y(n3061) );
 NOR2XLTS U1999 ( .A(n3067), .A(n3067_n), .B(n3068), .B(n3068_n), .Y(n3066_n), .Y(n3066) );
 NOR2XLTS U2000 ( .A(n2837), .A(n2837_n), .B(n2806), .B(n2806_n), .Y(n3067_n), .Y(n3067) );
 NOR2XLTS U2001 ( .A(n3098), .A(n3098_n), .B(n3099), .B(n3099_n), .Y(n3063_n), .Y(n3063) );
 NOR2XLTS U2002 ( .A(n3107), .A(n3107_n), .B(n3108), .B(n3108_n), .Y(n3106_n), .Y(n3106) );
 NOR2XLTS U2003 ( .A(n3109), .A(n3109_n), .B(n2781), .B(n2781_n), .Y(n3108_n), .Y(n3108) );
 NOR2XLTS U2004 ( .A(n3110), .A(n3110_n), .B(n2804), .B(n2804_n), .Y(n3107_n), .Y(n3107) );
 NOR2XLTS U2005 ( .A(n3111), .A(n3111_n), .B(n3112), .B(n3112_n), .Y(n3105_n), .Y(n3105) );
 NOR2XLTS U2006 ( .A(n2719), .A(n2719_n), .B(n2732), .B(n2732_n), .Y(n3111_n), .Y(n3111) );
 OR2XLTS U2007 ( .A(n2953), .A(n2953_n), .B(n3116), .B(n3116_n), .Y(n2963_n), .Y(n2963) );
 NOR2XLTS U2008 ( .A(n3119), .A(n3119_n), .B(n3120), .B(n3120_n), .Y(n3118_n), .Y(n3118) );
 NOR2XLTS U2009 ( .A(n3123), .A(n3123_n), .B(n3124), .B(n3124_n), .Y(n3122_n), .Y(n3122) );
 NOR2XLTS U2010 ( .A(n2705), .A(n2705_n), .B(n2790), .B(n2790_n), .Y(n3124_n), .Y(n3124) );
 NOR2XLTS U2011 ( .A(n3126), .A(n3126_n), .B(n3127), .B(n3127_n), .Y(n3121_n), .Y(n3121) );
 NOR2XLTS U2012 ( .A(n3133), .A(n3133_n), .B(n2735), .B(n2735_n), .Y(n3126_n), .Y(n3126) );
 NOR2XLTS U2013 ( .A(n2888), .A(n2888_n), .B(n3134), .B(n3134_n), .Y(n3133_n), .Y(n3133) );
 NOR2XLTS U2014 ( .A(n3135), .A(n3135_n), .B(n2815), .B(n2815_n), .Y(n3119_n), .Y(n3119) );
 NOR2XLTS U2015 ( .A(n3023), .A(n3023_n), .B(n3136), .B(n3136_n), .Y(n3135_n), .Y(n3135) );
 NOR2XLTS U2016 ( .A(n3137), .A(n3137_n), .B(n3138), .B(n3138_n), .Y(n3117_n), .Y(n3117) );
 NOR2XLTS U2017 ( .A(n2916), .A(n2916_n), .B(n2917), .B(n2917_n), .Y(n2915_n), .Y(n2915) );
 NOR2XLTS U2018 ( .A(n2997), .A(n2997_n), .B(n2998), .B(n2998_n), .Y(n2996_n), .Y(n2996) );
 NOR2XLTS U2019 ( .A(n3001), .A(n3001_n), .B(n3002), .B(n3002_n), .Y(n3000_n), .Y(n3000) );
 NOR2XLTS U2020 ( .A(n2977), .A(n2977_n), .B(n3003), .B(n3003_n), .Y(n3002_n), .Y(n3002) );
 NOR2XLTS U2021 ( .A(n3005), .A(n3005_n), .B(n2736), .B(n2736_n), .Y(n3001_n), .Y(n3001) );
 NOR2XLTS U2022 ( .A(n2881), .A(n2881_n), .B(n2748), .B(n2748_n), .Y(n3005_n), .Y(n3005) );
 NOR2XLTS U2023 ( .A(n3007), .A(n3007_n), .B(n3008), .B(n3008_n), .Y(n2999_n), .Y(n2999) );
 NOR2XLTS U2024 ( .A(n3011), .A(n3011_n), .B(n3012), .B(n3012_n), .Y(n3009_n), .Y(n3009) );
 NOR2XLTS U2025 ( .A(n2776), .A(n2776_n), .B(n2743), .B(n2743_n), .Y(n3012_n), .Y(n3012) );
 NOR2XLTS U2026 ( .A(n3014), .A(n3014_n), .B(n2801), .B(n2801_n), .Y(n3011_n), .Y(n3011) );
 NOR2XLTS U2027 ( .A(n3016), .A(n3016_n), .B(n2822), .B(n2822_n), .Y(n3007_n), .Y(n3007) );
 NOR2XLTS U2028 ( .A(n3019), .A(n3019_n), .B(n3020), .B(n3020_n), .Y(n2995_n), .Y(n2995) );
 NOR2XLTS U2029 ( .A(n3024), .A(n3024_n), .B(n3025), .B(n3025_n), .Y(n3021_n), .Y(n3021) );
 NOR2XLTS U2030 ( .A(n2759), .A(n2759_n), .B(n2771), .B(n2771_n), .Y(n3025_n), .Y(n3025) );
 NOR2XLTS U2031 ( .A(n2954), .A(n2954_n), .B(n2724), .B(n2724_n), .Y(n3024_n), .Y(n3024) );
 NOR2XLTS U2032 ( .A(n2920), .A(n2920_n), .B(n2921), .B(n2921_n), .Y(n2919_n), .Y(n2919) );
 NOR2XLTS U2033 ( .A(n2929), .A(n2929_n), .B(n2930), .B(n2930_n), .Y(n2918_n), .Y(n2918) );
 NOR2XLTS U2034 ( .A(n2942), .A(n2942_n), .B(n2943), .B(n2943_n), .Y(n2937_n), .Y(n2937) );
 NOR2XLTS U2035 ( .A(n2944), .A(n2944_n), .B(n2743), .B(n2743_n), .Y(n2943_n), .Y(n2943) );
 NOR2XLTS U2036 ( .A(n2763), .A(n2763_n), .B(n2848), .B(n2848_n), .Y(n2944_n), .Y(n2944) );
 NOR2XLTS U2037 ( .A(n2722), .A(n2722_n), .B(n2947), .B(n2947_n), .Y(n2942_n), .Y(n2942) );
 NOR2XLTS U2038 ( .A(n2948), .A(n2948_n), .B(n2949), .B(n2949_n), .Y(n2914_n), .Y(n2914) );
 NOR2XLTS U2039 ( .A(n3081), .A(n3081_n), .B(n3082), .B(n3082_n), .Y(n2951_n), .Y(n2951) );
 NOR2XLTS U2040 ( .A(n3086), .A(n3086_n), .B(n3087), .B(n3087_n), .Y(n3083_n), .Y(n3083) );
 NOR2XLTS U2041 ( .A(n3088), .A(n3088_n), .B(n2829), .B(n2829_n), .Y(n3086_n), .Y(n3086) );
 NOR2XLTS U2042 ( .A(n3093), .A(n3093_n), .B(n3094), .B(n3094_n), .Y(n3090_n), .Y(n3090) );
 NOR2XLTS U2043 ( .A(n3095), .A(n3095_n), .B(n2813), .B(n2813_n), .Y(n3094_n), .Y(n3094) );
 NOR2XLTS U2044 ( .A(n2778), .A(n2778_n), .B(n2869), .B(n2869_n), .Y(n3095_n), .Y(n3095) );
 NOR2XLTS U2045 ( .A(n3016), .A(n3016_n), .B(n2740), .B(n2740_n), .Y(n3093_n), .Y(n3093) );
 NOR2XLTS U2046 ( .A(n2816), .A(n2816_n), .B(n2784), .B(n2784_n), .Y(n3016_n), .Y(n3016) );
 NOR2XLTS U2047 ( .A(n2952), .A(n2952_n), .B(n2953), .B(n2953_n), .Y(n2950_n), .Y(n2950) );
 NOR2XLTS U2048 ( .A(n3146), .A(n3146_n), .B(n3147), .B(n3147_n), .Y(n3145_n), .Y(n3145) );
 NOR2XLTS U2049 ( .A(n3151), .A(n3151_n), .B(n2803), .B(n2803_n), .Y(n3146_n), .Y(n3146) );
 NOR2XLTS U2050 ( .A(n3152), .A(n3152_n), .B(n3153), .B(n3153_n), .Y(n3144_n), .Y(n3144) );
 NOR2XLTS U2051 ( .A(n2873), .A(n2873_n), .B(n2859), .B(n2859_n), .Y(n3158_n), .Y(n3158) );
 NOR2XLTS U2052 ( .A(n2750), .A(n2750_n), .B(n2863), .B(n2863_n), .Y(n2982_n), .Y(n2982) );
 NOR2XLTS U2053 ( .A(n2838), .A(n2838_n), .B(n2802), .B(n2802_n), .Y(n2952_n), .Y(n2952) );
 NOR2XLTS U2054 ( .A(n2957), .A(n2957_n), .B(n2958), .B(n2958_n), .Y(n2956_n), .Y(n2956) );
 NOR2XLTS U2055 ( .A(n3071), .A(n3071_n), .B(n3072), .B(n3072_n), .Y(n2959_n), .Y(n2959) );
 NOR2XLTS U2056 ( .A(n3078), .A(n3078_n), .B(n3079), .B(n3079_n), .Y(n3075_n), .Y(n3075) );
 NOR2XLTS U2057 ( .A(n2715), .A(n2715_n), .B(n2776), .B(n2776_n), .Y(n3079_n), .Y(n3079) );
 NOR2XLTS U2058 ( .A(n2757), .A(n2757_n), .B(n2826), .B(n2826_n), .Y(n3078_n), .Y(n3078) );
 NOR2XLTS U2059 ( .A(n3247), .A(n3247_n), .B(n3508), .B(n3508_n), .Y(n3164_n), .Y(n3164) );
 OR2XLTS U2060 ( .A(n3057), .A(n3057_n), .B(n3509), .B(n3509_n), .Y(n3508_n), .Y(n3508) );
 NOR2XLTS U2061 ( .A(n3512), .A(n3512_n), .B(n3513), .B(n3513_n), .Y(n3511_n), .Y(n3511) );
 NOR2XLTS U2062 ( .A(n3516), .A(n3516_n), .B(n3517), .B(n3517_n), .Y(n3514_n), .Y(n3514) );
 NOR2XLTS U2063 ( .A(n3187), .A(n3187_n), .B(n2772), .B(n2772_n), .Y(n3517_n), .Y(n3517) );
 NOR2XLTS U2064 ( .A(n3518), .A(n3518_n), .B(n2768), .B(n2768_n), .Y(n3516_n), .Y(n3516) );
 NOR2XLTS U2065 ( .A(n2842), .A(n2842_n), .B(n2786), .B(n2786_n), .Y(n3518_n), .Y(n3518) );
 NOR2XLTS U2066 ( .A(n3218), .A(n3218_n), .B(n2752), .B(n2752_n), .Y(n3512_n), .Y(n3512) );
 NOR2XLTS U2067 ( .A(n3519), .A(n3519_n), .B(n3520), .B(n3520_n), .Y(n3510_n), .Y(n3510) );
 INVXLTS U2068 ( .A(n3222), .A(n3222_n), .Y(n3458_n), .Y(n3458) );
 NOR2XLTS U2069 ( .A(n3525), .A(n3525_n), .B(n2828), .B(n2828_n), .Y(n3519_n), .Y(n3519) );
 NOR2XLTS U2070 ( .A(n2702), .A(n2702_n), .B(n3136), .B(n3136_n), .Y(n3525_n), .Y(n3525) );
 NOR2XLTS U2071 ( .A(n3530), .A(n3530_n), .B(n3531), .B(n3531_n), .Y(n3529_n), .Y(n3529) );
 NOR2XLTS U2072 ( .A(n3151), .A(n3151_n), .B(n2736), .B(n2736_n), .Y(n3531_n), .Y(n3531) );
 NOR2XLTS U2073 ( .A(n3532), .A(n3532_n), .B(n2732), .B(n2732_n), .Y(n3530_n), .Y(n3530) );
 NOR2XLTS U2074 ( .A(n2875), .A(n2875_n), .B(n3424), .B(n3424_n), .Y(n3532_n), .Y(n3532) );
 NOR2XLTS U2075 ( .A(n3533), .A(n3533_n), .B(n3534), .B(n3534_n), .Y(n3528_n), .Y(n3528) );
 NOR2XLTS U2076 ( .A(n3536), .A(n3536_n), .B(n3537), .B(n3537_n), .Y(n3535_n), .Y(n3535) );
 NOR2XLTS U2077 ( .A(n2704), .A(n2704_n), .B(n2802), .B(n2802_n), .Y(n3537_n), .Y(n3537) );
 NOR2XLTS U2078 ( .A(n3169), .A(n3169_n), .B(n2834), .B(n2834_n), .Y(n3536_n), .Y(n3536) );
 NOR2XLTS U2079 ( .A(n3110), .A(n3110_n), .B(n2807), .B(n2807_n), .Y(n3533_n), .Y(n3533) );
 INVXLTS U2080 ( .A(n3136), .A(n3136_n), .Y(n3110_n), .Y(n3110) );
 NOR2XLTS U2081 ( .A(n2740), .A(n2740_n), .B(n2723), .B(n2723_n), .Y(n3172_n), .Y(n3172) );
 NOR2XLTS U2082 ( .A(n3175), .A(n3175_n), .B(n3176), .B(n3176_n), .Y(n3174_n), .Y(n3174) );
 NOR2XLTS U2083 ( .A(n3432), .A(n3432_n), .B(n3433), .B(n3433_n), .Y(n3430_n), .Y(n3430) );
 NOR2XLTS U2084 ( .A(n3179), .A(n3179_n), .B(n3180), .B(n3180_n), .Y(n3178_n), .Y(n3178) );
 INVXLTS U2085 ( .A(n3184), .A(n3184_n), .Y(n3183_n), .Y(n3183) );
 NOR2XLTS U2086 ( .A(n3185), .A(n3185_n), .B(n3186), .B(n3186_n), .Y(n3181_n), .Y(n3181) );
 NOR2XLTS U2087 ( .A(n3187), .A(n3187_n), .B(n2826), .B(n2826_n), .Y(n3186_n), .Y(n3186) );
 NOR2XLTS U2088 ( .A(n2873), .A(n2873_n), .B(n2877), .B(n2877_n), .Y(n3187_n), .Y(n3187) );
 NOR2XLTS U2089 ( .A(n3188), .A(n3188_n), .B(n2813), .B(n2813_n), .Y(n3185_n), .Y(n3185) );
 NOR2XLTS U2090 ( .A(n2887), .A(n2887_n), .B(n2879), .B(n2879_n), .Y(n3188_n), .Y(n3188) );
 NOR2XLTS U2091 ( .A(n3189), .A(n3189_n), .B(n3190), .B(n3190_n), .Y(n3177_n), .Y(n3177) );
 NOR2XLTS U2092 ( .A(n3195), .A(n3195_n), .B(n2705), .B(n2705_n), .Y(n3189_n), .Y(n3189) );
 NOR2XLTS U2093 ( .A(n2845), .A(n2845_n), .B(n2934), .B(n2934_n), .Y(n3195_n), .Y(n3195) );
 NOR2XLTS U2094 ( .A(n3196), .A(n3196_n), .B(n3197), .B(n3197_n), .Y(n3173_n), .Y(n3173) );
 NOR2XLTS U2095 ( .A(n3200), .A(n3200_n), .B(n3201), .B(n3201_n), .Y(n3198_n), .Y(n3198) );
 NOR2XLTS U2096 ( .A(n2819), .A(n2819_n), .B(n2835), .B(n2835_n), .Y(n3201_n), .Y(n3201) );
 NOR2XLTS U2097 ( .A(n2801), .A(n2801_n), .B(n2752), .B(n2752_n), .Y(n3200_n), .Y(n3200) );
 NOR2XLTS U2098 ( .A(n3087), .A(n3087_n), .B(n3206), .B(n3206_n), .Y(n3205_n), .Y(n3205) );
 NOR2XLTS U2099 ( .A(n2830), .A(n2830_n), .B(n2742), .B(n2742_n), .Y(n3206_n), .Y(n3206) );
 NOR2XLTS U2100 ( .A(n2760), .A(n2760_n), .B(n2721), .B(n2721_n), .Y(n3087_n), .Y(n3087) );
 NOR2XLTS U2101 ( .A(n3207), .A(n3207_n), .B(n3208), .B(n3208_n), .Y(n3204_n), .Y(n3204) );
 NOR2XLTS U2102 ( .A(n3015), .A(n3015_n), .B(n2827), .B(n2827_n), .Y(n3208_n), .Y(n3208) );
 NOR2XLTS U2103 ( .A(n3104), .A(n3104_n), .B(n2789), .B(n2789_n), .Y(n3207_n), .Y(n3207) );
 NOR2XLTS U2104 ( .A(n3211), .A(n3211_n), .B(n3212), .B(n3212_n), .Y(n3210_n), .Y(n3210) );
 NOR2XLTS U2105 ( .A(n3184), .A(n3184_n), .B(n2835), .B(n2835_n), .Y(n3212_n), .Y(n3212) );
 NOR2XLTS U2106 ( .A(n2764), .A(n2764_n), .B(n2841), .B(n2841_n), .Y(n3184_n), .Y(n3184) );
 NOR2XLTS U2107 ( .A(n3213), .A(n3213_n), .B(n2795), .B(n2795_n), .Y(n3211_n), .Y(n3211) );
 NOR2XLTS U2108 ( .A(n2933), .A(n2933_n), .B(n3166), .B(n3166_n), .Y(n3213_n), .Y(n3213) );
 NOR2XLTS U2109 ( .A(n3214), .A(n3214_n), .B(n3215), .B(n3215_n), .Y(n3209_n), .Y(n3209) );
 NOR2XLTS U2110 ( .A(n3218), .A(n3218_n), .B(n2807), .B(n2807_n), .Y(n3214_n), .Y(n3214) );
 NOR2XLTS U2111 ( .A(n2779), .A(n2779_n), .B(n2882), .B(n2882_n), .Y(n3218_n), .Y(n3218) );
 NOR2XLTS U2112 ( .A(n3364), .A(n3364_n), .B(n3489), .B(n3489_n), .Y(n3488_n), .Y(n3488) );
 NOR2XLTS U2113 ( .A(n3492), .A(n3492_n), .B(n3493), .B(n3493_n), .Y(n3490_n), .Y(n3490) );
 NOR2XLTS U2114 ( .A(n2829), .A(n2829_n), .B(n2722), .B(n2722_n), .Y(n3493_n), .Y(n3493) );
 NOR2XLTS U2115 ( .A(n2780), .A(n2780_n), .B(n2792), .B(n2792_n), .Y(n3492_n), .Y(n3492) );
 NOR2XLTS U2116 ( .A(n3494), .A(n3494_n), .B(n3495), .B(n3495_n), .Y(n3487_n), .Y(n3487) );
 NOR2XLTS U2117 ( .A(n2717), .A(n2717_n), .B(n2756), .B(n2756_n), .Y(n3498_n), .Y(n3498) );
 NOR2XLTS U2118 ( .A(n2769), .A(n2769_n), .B(n2849), .B(n2849_n), .Y(n3047_n), .Y(n3047) );
 NOR2XLTS U2119 ( .A(n3504), .A(n3504_n), .B(n3505), .B(n3505_n), .Y(n3501_n), .Y(n3501) );
 NOR2XLTS U2120 ( .A(n3506), .A(n3506_n), .B(n2753), .B(n2753_n), .Y(n3505_n), .Y(n3505) );
 NOR2XLTS U2121 ( .A(n2878), .A(n2878_n), .B(n2744), .B(n2744_n), .Y(n3506_n), .Y(n3506) );
 NOR2XLTS U2122 ( .A(n3507), .A(n3507_n), .B(n2724), .B(n2724_n), .Y(n3504_n), .Y(n3504) );
 NOR2XLTS U2123 ( .A(n2883), .A(n2883_n), .B(n2725), .B(n2725_n), .Y(n3507_n), .Y(n3507) );
 NOR2XLTS U2124 ( .A(n3225), .A(n3225_n), .B(n2715), .B(n2715_n), .Y(n3224_n), .Y(n3224) );
 NOR2XLTS U2125 ( .A(n2809), .A(n2809_n), .B(n2934), .B(n2934_n), .Y(n3225_n), .Y(n3225) );
 NOR2XLTS U2126 ( .A(n2813), .A(n2813_n), .B(n3167), .B(n3167_n), .Y(n3223_n), .Y(n3223) );
 NOR2XLTS U2127 ( .A(n3226), .A(n3226_n), .B(n3227), .B(n3227_n), .Y(n3031_n), .Y(n3031) );
 NOR2XLTS U2128 ( .A(n3230), .A(n3230_n), .B(n3231), .B(n3231_n), .Y(n3228_n), .Y(n3228) );
 NOR2XLTS U2129 ( .A(n2881), .A(n2881_n), .B(n2860), .B(n2860_n), .Y(n3088_n), .Y(n3088) );
 NOR2XLTS U2130 ( .A(n3235), .A(n3235_n), .B(n2796), .B(n2796_n), .Y(n3230_n), .Y(n3230) );
 NOR2XLTS U2131 ( .A(n2879), .A(n2879_n), .B(n2747), .B(n2747_n), .Y(n3235_n), .Y(n3235) );
 NOR2XLTS U2132 ( .A(n3238), .A(n3238_n), .B(n3239), .B(n3239_n), .Y(n3237_n), .Y(n3237) );
 AND2XLTS U2133 ( .A(n3244), .A(n3244_n), .B(n3245), .B(n3245_n), .Y(n3242_n), .Y(n3242) );
 INVXLTS U2134 ( .A(n2839), .A(n2839_n), .Y(n3004_n), .Y(n3004) );
 NOR2XLTS U2135 ( .A(n3123), .A(n3123_n), .B(n3246), .B(n3246_n), .Y(n3236_n), .Y(n3236) );
 NOR2XLTS U2136 ( .A(n3109), .A(n3109_n), .B(n2734), .B(n2734_n), .Y(n3246_n), .Y(n3246) );
 NOR2XLTS U2137 ( .A(n3202), .A(n3202_n), .B(n2828), .B(n2828_n), .Y(n3123_n), .Y(n3123) );
 NOR2XLTS U2138 ( .A(n3438), .A(n3438_n), .B(n3439), .B(n3439_n), .Y(n3248_n), .Y(n3248) );
 OR2XLTS U2139 ( .A(n3440), .A(n3440_n), .B(n3441), .B(n3441_n), .Y(n3439_n), .Y(n3439) );
 NOR2XLTS U2140 ( .A(n3450), .A(n3450_n), .B(n3451), .B(n3451_n), .Y(n3449_n), .Y(n3449) );
 NOR2XLTS U2141 ( .A(n3222), .A(n3222_n), .B(n2733), .B(n2733_n), .Y(n3451_n), .Y(n3451) );
 NOR2XLTS U2142 ( .A(n3171), .A(n3171_n), .B(n2793), .B(n2793_n), .Y(n3450_n), .Y(n3450) );
 NOR2XLTS U2143 ( .A(n3452), .A(n3452_n), .B(n3453), .B(n3453_n), .Y(n3448_n), .Y(n3448) );
 NOR2XLTS U2144 ( .A(n3456), .A(n3456_n), .B(n3457), .B(n3457_n), .Y(n3454_n), .Y(n3454) );
 NOR2XLTS U2145 ( .A(n2796), .A(n2796_n), .B(n2835), .B(n2835_n), .Y(n3457_n), .Y(n3457) );
 NOR2XLTS U2146 ( .A(n2767), .A(n2767_n), .B(n2814), .B(n2814_n), .Y(n3456_n), .Y(n3456) );
 NOR2XLTS U2147 ( .A(n2941), .A(n2941_n), .B(n2824), .B(n2824_n), .Y(n3452_n), .Y(n3452) );
 NOR2XLTS U2148 ( .A(n2852), .A(n2852_n), .B(n2855), .B(n2855_n), .Y(n2941_n), .Y(n2941) );
 NOR2XLTS U2149 ( .A(n3251), .A(n3251_n), .B(n3252), .B(n3252_n), .Y(n3250_n), .Y(n3250) );
 NOR2XLTS U2150 ( .A(n3259), .A(n3259_n), .B(n3260), .B(n3260_n), .Y(n3249_n), .Y(n3249) );
 NOR2XLTS U2151 ( .A(n3059), .A(n3059_n), .B(n3540), .B(n3540_n), .Y(n3539_n), .Y(n3539) );
 NOR2XLTS U2152 ( .A(n3545), .A(n3545_n), .B(n3546), .B(n3546_n), .Y(n3541_n), .Y(n3541) );
 INVXLTS U2153 ( .A(n3134), .A(n3134_n), .Y(n3040_n), .Y(n3040) );
 NOR2XLTS U2154 ( .A(n2873), .A(n2873_n), .B(n2779), .B(n2779_n), .Y(n3544_n), .Y(n3544) );
 NOR2XLTS U2155 ( .A(n3564), .A(n3564_n), .B(n3565), .B(n3565_n), .Y(n3557_n), .Y(n3557) );
 NOR2XLTS U2156 ( .A(n3572), .A(n3572_n), .B(n2757), .B(n2757_n), .Y(n3564_n), .Y(n3564) );
 NOR2XLTS U2157 ( .A(n2810), .A(n2810_n), .B(n3574), .B(n3574_n), .Y(n3572_n), .Y(n3572) );
 NOR2XLTS U2158 ( .A(n3058), .A(n3058_n), .B(n3575), .B(n3575_n), .Y(n3538_n), .Y(n3538) );
 NOR2XLTS U2159 ( .A(n3411), .A(n3411_n), .B(n3582), .B(n3582_n), .Y(n3581_n), .Y(n3581) );
 NOR2XLTS U2160 ( .A(n2822), .A(n2822_n), .B(n2771), .B(n2771_n), .Y(n3582_n), .Y(n3582) );
 NOR2XLTS U2161 ( .A(n3584), .A(n3584_n), .B(n3585), .B(n3585_n), .Y(n3580_n), .Y(n3580) );
 NOR2XLTS U2162 ( .A(n3171), .A(n3171_n), .B(n2805), .B(n2805_n), .Y(n3585_n), .Y(n3585) );
 NOR2XLTS U2163 ( .A(n2858), .A(n2858_n), .B(n2745), .B(n2745_n), .Y(n3171_n), .Y(n3171) );
 NOR2XLTS U2164 ( .A(n3588), .A(n3588_n), .B(n2720), .B(n2720_n), .Y(n3584_n), .Y(n3584) );
 NOR2XLTS U2165 ( .A(n2817), .A(n2817_n), .B(n2854), .B(n2854_n), .Y(n3588_n), .Y(n3588) );
 NOR2XLTS U2166 ( .A(n3270), .A(n3270_n), .B(n3271), .B(n3271_n), .Y(n3269_n), .Y(n3269) );
 NOR2XLTS U2167 ( .A(n2957), .A(n2957_n), .B(n2968), .B(n2968_n), .Y(n3273_n), .Y(n3273) );
 NOR2XLTS U2168 ( .A(n3276), .A(n3276_n), .B(n3277), .B(n3277_n), .Y(n3275_n), .Y(n3275) );
 NOR2XLTS U2169 ( .A(n3282), .A(n3282_n), .B(n3036), .B(n3036_n), .Y(n3280_n), .Y(n3280) );
 NOR2XLTS U2170 ( .A(n2800), .A(n2800_n), .B(n2814), .B(n2814_n), .Y(n3036_n), .Y(n3036) );
 NOR2XLTS U2171 ( .A(n2826), .A(n2826_n), .B(n2742), .B(n2742_n), .Y(n3282_n), .Y(n3282) );
 NOR2XLTS U2172 ( .A(n3283), .A(n3283_n), .B(n3284), .B(n3284_n), .Y(n3274_n), .Y(n3274) );
 INVXLTS U2173 ( .A(n3288), .A(n3288_n), .Y(n3104_n), .Y(n3104) );
 NOR2XLTS U2174 ( .A(n2912), .A(n2912_n), .B(n3289), .B(n3289_n), .Y(n3132_n), .Y(n3132) );
 NOR2XLTS U2175 ( .A(n3293), .A(n3293_n), .B(n3294), .B(n3294_n), .Y(n3290_n), .Y(n3290) );
 NOR2XLTS U2176 ( .A(n3109), .A(n3109_n), .B(n2766), .B(n2766_n), .Y(n3294_n), .Y(n3294) );
 NOR2XLTS U2177 ( .A(n2717), .A(n2717_n), .B(n2738), .B(n2738_n), .Y(n3109_n), .Y(n3109) );
 NOR2XLTS U2178 ( .A(n3295), .A(n3295_n), .B(n2861), .B(n2861_n), .Y(n3293_n), .Y(n3293) );
 NOR2XLTS U2179 ( .A(n3298), .A(n3298_n), .B(n3299), .B(n3299_n), .Y(n3297_n), .Y(n3297) );
 NOR2XLTS U2180 ( .A(n2954), .A(n2954_n), .B(n2831), .B(n2831_n), .Y(n3299_n), .Y(n3299) );
 NOR2XLTS U2181 ( .A(n2806), .A(n2806_n), .B(n2822), .B(n2822_n), .Y(n3298_n), .Y(n3298) );
 NOR2XLTS U2182 ( .A(n3300), .A(n3300_n), .B(n3301), .B(n3301_n), .Y(n3296_n), .Y(n3296) );
 NOR2XLTS U2183 ( .A(n2794), .A(n2794_n), .B(n2710), .B(n2710_n), .Y(n3300_n), .Y(n3300) );
 NOR2XLTS U2184 ( .A(n3305), .A(n3305_n), .B(n3306), .B(n3306_n), .Y(n3272_n), .Y(n3272) );
 NOR2XLTS U2185 ( .A(n3309), .A(n3309_n), .B(n3310), .B(n3310_n), .Y(n3308_n), .Y(n3308) );
 NOR2XLTS U2186 ( .A(n2716), .A(n2716_n), .B(n2805), .B(n2805_n), .Y(n3310_n), .Y(n3310) );
 NOR2XLTS U2187 ( .A(n2710), .A(n2710_n), .B(n2827), .B(n2827_n), .Y(n3309_n), .Y(n3309) );
 NOR2XLTS U2188 ( .A(n3311), .A(n3311_n), .B(n3312), .B(n3312_n), .Y(n3307_n), .Y(n3307) );
 NOR2XLTS U2189 ( .A(n2720), .A(n2720_n), .B(n2815), .B(n2815_n), .Y(n3312_n), .Y(n3312) );
 NOR2XLTS U2190 ( .A(n3151), .A(n3151_n), .B(n2775), .B(n2775_n), .Y(n3311_n), .Y(n3311) );
 NOR2XLTS U2191 ( .A(n2730), .A(n2730_n), .B(n3085), .B(n3085_n), .Y(n3151_n), .Y(n3151) );
 NOR2XLTS U2192 ( .A(n3315), .A(n3315_n), .B(n3316), .B(n3316_n), .Y(n3314_n), .Y(n3314) );
 NOR2XLTS U2193 ( .A(n3014), .A(n3014_n), .B(n2833), .B(n2833_n), .Y(n3316_n), .Y(n3316) );
 NOR2XLTS U2194 ( .A(n2693), .A(n2693_n), .B(n2765), .B(n2765_n), .Y(n3014_n), .Y(n3014) );
 NOR2XLTS U2195 ( .A(n3317), .A(n3317_n), .B(n2790), .B(n2790_n), .Y(n3315_n), .Y(n3315) );
 NOR2XLTS U2196 ( .A(n2701), .A(n2701_n), .B(n3257), .B(n3257_n), .Y(n3317_n), .Y(n3317) );
 NOR2XLTS U2197 ( .A(n3318), .A(n3318_n), .B(n3319), .B(n3319_n), .Y(n3313_n), .Y(n3313) );
 NOR2XLTS U2198 ( .A(n3320), .A(n3320_n), .B(n2727), .B(n2727_n), .Y(n3319_n), .Y(n3319) );
 NOR2XLTS U2199 ( .A(n2844), .A(n2844_n), .B(n2851), .B(n2851_n), .Y(n3320_n), .Y(n3320) );
 NOR2XLTS U2200 ( .A(n3321), .A(n3321_n), .B(n2800), .B(n2800_n), .Y(n3318_n), .Y(n3318) );
 NOR2XLTS U2201 ( .A(n2783), .A(n2783_n), .B(n2809), .B(n2809_n), .Y(n3321_n), .Y(n3321) );
 OR2XLTS U2202 ( .A(n3019), .A(n3019_n), .B(n3322), .B(n3322_n), .Y(n3270_n), .Y(n3270) );
 NOR2XLTS U2203 ( .A(n3324), .A(n3324_n), .B(n3325), .B(n3325_n), .Y(n3323_n), .Y(n3323) );
 NOR2XLTS U2204 ( .A(n2762), .A(n2762_n), .B(n2742), .B(n2742_n), .Y(n3325_n), .Y(n3325) );
 NOR2XLTS U2205 ( .A(n2820), .A(n2820_n), .B(n2759), .B(n2759_n), .Y(n3324_n), .Y(n3324) );
 NOR2XLTS U2206 ( .A(n3326), .A(n3326_n), .B(n3327), .B(n3327_n), .Y(n2960_n), .Y(n2960) );
 NOR2XLTS U2207 ( .A(n2798), .A(n2798_n), .B(n2738), .B(n2738_n), .Y(n2977_n), .Y(n2977) );
 NOR2XLTS U2208 ( .A(n3334), .A(n3334_n), .B(n3335), .B(n3335_n), .Y(n3331_n), .Y(n3331) );
 NOR2XLTS U2209 ( .A(n3336), .A(n3336_n), .B(n2793), .B(n2793_n), .Y(n3335_n), .Y(n3335) );
 NOR2XLTS U2210 ( .A(n2882), .A(n2882_n), .B(n2870), .B(n2870_n), .Y(n3336_n), .Y(n3336) );
 NOR2XLTS U2211 ( .A(n3337), .A(n3337_n), .B(n2834), .B(n2834_n), .Y(n3334_n), .Y(n3334) );
 NOR2XLTS U2212 ( .A(n2718), .A(n2718_n), .B(n2816), .B(n2816_n), .Y(n3337_n), .Y(n3337) );
 NOR2XLTS U2213 ( .A(n3340), .A(n3340_n), .B(n3341), .B(n3341_n), .Y(n3339_n), .Y(n3339) );
 INVXLTS U2214 ( .A(n2740), .A(n2740_n), .Y(n3023_n), .Y(n3023) );
 NOR2XLTS U2215 ( .A(n3345), .A(n3345_n), .B(n3346), .B(n3346_n), .Y(n3338_n), .Y(n3338) );
 NOR2XLTS U2216 ( .A(n2871), .A(n2871_n), .B(n2859), .B(n2859_n), .Y(n3350_n), .Y(n3350) );
 NOR2XLTS U2217 ( .A(n2695), .A(n2695_n), .B(n2713), .B(n2713_n), .Y(n3169_n), .Y(n3169) );
 INVXLTS U2218 ( .A(n2792), .A(n2792_n), .Y(n3097_n), .Y(n3097) );
 INVXLTS U2219 ( .A(n2795), .A(n2795_n), .Y(n2924_n), .Y(n2924) );
 NOR2XLTS U2220 ( .A(n2797), .A(n2797_n), .B(n2842), .B(n2842_n), .Y(n3295_n), .Y(n3295) );
 NOR2XLTS U2221 ( .A(n3523), .A(n3523_n), .B(n3289), .B(n3289_n), .Y(n2986_n), .Y(n2986) );
 NOR2XLTS U2222 ( .A(n2811), .A(n2811_n), .B(n2714), .B(n2714_n), .Y(n3222_n), .Y(n3222) );
 NOR2XLTS U2223 ( .A(n3568), .A(n3568_n), .B(n3573), .B(n3573_n), .Y(n2928_n), .Y(n2928) );
 NOR2XLTS U2224 ( .A(n3363), .A(n3363_n), .B(n2788), .B(n2788_n), .Y(n3357_n), .Y(n3357) );
 NOR2XLTS U2225 ( .A(n2869), .A(n2869_n), .B(n2696), .B(n2696_n), .Y(n3363_n), .Y(n3363) );
 INVXLTS U2226 ( .A(n2824), .A(n2824_n), .Y(n3006_n), .Y(n3006) );
 NOR2XLTS U2227 ( .A(n3364), .A(n3364_n), .B(n3365), .B(n3365_n), .Y(n3017_n), .Y(n3017) );
 NOR2XLTS U2228 ( .A(n3368), .A(n3368_n), .B(n3369), .B(n3369_n), .Y(n3366_n), .Y(n3366) );
 NOR2XLTS U2229 ( .A(n2830), .A(n2830_n), .B(n2710), .B(n2710_n), .Y(n3369_n), .Y(n3369) );
 NOR2XLTS U2230 ( .A(n2803), .A(n2803_n), .B(n3167), .B(n3167_n), .Y(n3368_n), .Y(n3368) );
 NOR2XLTS U2231 ( .A(n2821), .A(n2821_n), .B(n2823), .B(n2823_n), .Y(n3364_n), .Y(n3364) );
 NOR2XLTS U2232 ( .A(n3371), .A(n3371_n), .B(n3372), .B(n3372_n), .Y(n2955_n), .Y(n2955) );
 NOR2XLTS U2233 ( .A(n3375), .A(n3375_n), .B(n3376), .B(n3376_n), .Y(n3374_n), .Y(n3374) );
 NOR2XLTS U2234 ( .A(n2835), .A(n2835_n), .B(n2731), .B(n2731_n), .Y(n3376_n), .Y(n3376) );
 NOR2XLTS U2235 ( .A(n2739), .A(n2739_n), .B(n2752), .B(n2752_n), .Y(n3375_n), .Y(n3375) );
 NOR2XLTS U2236 ( .A(n3377), .A(n3377_n), .B(n3378), .B(n3378_n), .Y(n3373_n), .Y(n3373) );
 NOR2XLTS U2237 ( .A(n2733), .A(n2733_n), .B(n2789), .B(n2789_n), .Y(n3377_n), .Y(n3377) );
 NOR2XLTS U2238 ( .A(n3382), .A(n3382_n), .B(n3383), .B(n3383_n), .Y(n3381_n), .Y(n3381) );
 NOR2XLTS U2239 ( .A(n2711), .A(n2711_n), .B(n2762), .B(n2762_n), .Y(n3383_n), .Y(n3383) );
 NOR2XLTS U2240 ( .A(n3384), .A(n3384_n), .B(n2791), .B(n2791_n), .Y(n3382_n), .Y(n3382) );
 NOR2XLTS U2241 ( .A(n2886), .A(n2886_n), .B(n2862), .B(n2862_n), .Y(n3384_n), .Y(n3384) );
 NOR2XLTS U2242 ( .A(n3385), .A(n3385_n), .B(n3386), .B(n3386_n), .Y(n3380_n), .Y(n3380) );
 NOR2XLTS U2243 ( .A(n3390), .A(n3390_n), .B(n2820), .B(n2820_n), .Y(n3385_n), .Y(n3385) );
 NOR2XLTS U2244 ( .A(n2729), .A(n2729_n), .B(n3115), .B(n3115_n), .Y(n3390_n), .Y(n3390) );
 NOR2XLTS U2245 ( .A(n3392), .A(n3392_n), .B(n3393), .B(n3393_n), .Y(n3018_n), .Y(n3018) );
 NOR2XLTS U2246 ( .A(n2909), .A(n2909_n), .B(n2912), .B(n2912_n), .Y(n3561_n), .Y(n3561) );
 INVXLTS U2247 ( .A(n2734), .A(n2734_n), .Y(n3085_n), .Y(n3085) );
 NOR2XLTS U2248 ( .A(n3402), .A(n3402_n), .B(n3403), .B(n3403_n), .Y(n3399_n), .Y(n3399) );
 NOR2XLTS U2249 ( .A(n3404), .A(n3404_n), .B(n2761), .B(n2761_n), .Y(n3403_n), .Y(n3403) );
 NOR2XLTS U2250 ( .A(n3405), .A(n3405_n), .B(n2728), .B(n2728_n), .Y(n3402_n), .Y(n3402) );
 NOR2XLTS U2251 ( .A(n2841), .A(n2841_n), .B(n2737), .B(n2737_n), .Y(n3405_n), .Y(n3405) );
 NOR2XLTS U2252 ( .A(n3406), .A(n3406_n), .B(n3407), .B(n3407_n), .Y(n2965_n), .Y(n2965) );
 NOR2XLTS U2253 ( .A(n3410), .A(n3410_n), .B(n3411), .B(n3411_n), .Y(n3409_n), .Y(n3409) );
 NOR2XLTS U2254 ( .A(n2802), .A(n2802_n), .B(n2834), .B(n2834_n), .Y(n3411_n), .Y(n3411) );
 NOR2XLTS U2255 ( .A(n2723), .A(n2723_n), .B(n2733), .B(n2733_n), .Y(n3410_n), .Y(n3410) );
 NOR2XLTS U2256 ( .A(n3412), .A(n3412_n), .B(n3413), .B(n3413_n), .Y(n3408_n), .Y(n3408) );
 NOR2XLTS U2257 ( .A(n2731), .A(n2731_n), .B(n2823), .B(n2823_n), .Y(n3413_n), .Y(n3413) );
 INVXLTS U2258 ( .A(n3398), .A(n3398_n), .Y(n3304_n), .Y(n3304) );
 NOR2XLTS U2259 ( .A(n2727), .A(n2727_n), .B(n2814), .B(n2814_n), .Y(n3412_n), .Y(n3412) );
 NOR2XLTS U2260 ( .A(n3416), .A(n3416_n), .B(n3417), .B(n3417_n), .Y(n3415_n), .Y(n3415) );
 NOR2XLTS U2261 ( .A(n3418), .A(n3418_n), .B(n2772), .B(n2772_n), .Y(n3417_n), .Y(n3417) );
 NOR2XLTS U2262 ( .A(n3461), .A(n3461_n), .B(n3583), .B(n3583_n), .Y(n3051_n), .Y(n3051) );
 INVXLTS U2263 ( .A(n3499), .A(n3499_n), .Y(n3461_n), .Y(n3461) );
 NOR2XLTS U2264 ( .A(n2857), .A(n2857_n), .B(n3288), .B(n3288_n), .Y(n3418_n), .Y(n3418) );
 NOR2XLTS U2265 ( .A(n3523), .A(n3523_n), .B(n3524), .B(n3524_n), .Y(n2975_n), .Y(n2975) );
 NOR2XLTS U2266 ( .A(n3556), .A(n3556_n), .B(n3289), .B(n3289_n), .Y(n2939_n), .Y(n2939) );
 NOR2XLTS U2267 ( .A(n3419), .A(n3419_n), .B(n2806), .B(n2806_n), .Y(n3416_n), .Y(n3416) );
 NOR2XLTS U2268 ( .A(n2903), .A(n2903_n), .B(n3398), .B(n3398_n), .Y(n2946_n), .Y(n2946) );
 NOR2XLTS U2269 ( .A(n2874), .A(n2874_n), .B(n2862), .B(n2862_n), .Y(n3419_n), .Y(n3419) );
 NOR2XLTS U2270 ( .A(n3526), .A(n3526_n), .B(n3527), .B(n3527_n), .Y(n2933_n), .Y(n2933) );
 NOR2XLTS U2271 ( .A(n3523), .A(n3523_n), .B(n3563), .B(n3563_n), .Y(n2994_n), .Y(n2994) );
 OR2XLTS U2272 ( .A(n2891), .A(n2891_n), .B(n2908), .B(n2908_n), .Y(n3563_n), .Y(n3563) );
 INVXLTS U2273 ( .A(n3466), .A(n3466_n), .Y(n3523_n), .Y(n3523) );
 NOR2XLTS U2274 ( .A(n3420), .A(n3420_n), .B(n3421), .B(n3421_n), .Y(n3414_n), .Y(n3414) );
 NOR2XLTS U2275 ( .A(n3556), .A(n3556_n), .B(n3524), .B(n3524_n), .Y(n2925_n), .Y(n2925) );
 NOR2XLTS U2276 ( .A(n3526), .A(n3526_n), .B(n3556), .B(n3556_n), .Y(n3077_n), .Y(n3077) );
 INVXLTS U2277 ( .A(n2729), .A(n2729_n), .Y(n3015_n), .Y(n3015) );
 NOR2XLTS U2278 ( .A(n2708), .A(n2708_n), .B(n3583), .B(n3583_n), .Y(n3161_n), .Y(n3161) );
 INVXLTS U2279 ( .A(n3586), .A(n3586_n), .Y(n3583_n), .Y(n3583) );
 NOR2XLTS U2280 ( .A(n2893), .A(n2893_n), .B(n2906), .B(n2906_n), .Y(n3586_n), .Y(n3586) );
 NOR2XLTS U2281 ( .A(n3426), .A(n3426_n), .B(n3427), .B(n3427_n), .Y(n3420_n), .Y(n3420) );
 AND2XLTS U2282 ( .A(n2899), .A(n2899_n), .B(n2902), .B(n2902_n), .Y(n3428_n), .Y(n3428) );
 NOR2XLTS U2283 ( .A(n2911), .A(n2911_n), .B(n3570), .B(n3570_n), .Y(n3587_n), .Y(n3587) );
 INVXLTS U2284 ( .A(n3568), .A(n3568_n), .Y(n3560_n), .Y(n3560) );
 OR2XLTS U2285 ( .A(n2896), .A(n2896_n), .B(n2891), .B(n2891_n), .Y(n3568_n), .Y(n3568) );
 NOR2XLTS U2286 ( .A(n2896), .A(n2896_n), .B(n3289), .B(n3289_n), .Y(n3446_n), .Y(n3446) );
 INVXLTS U2287 ( .A(n2908), .A(n2908_n), .Y(n3570_n), .Y(n3570) );
 NOR2XLTS U2288 ( .A(n3526), .A(n3526_n), .B(n3578), .B(n3578_n), .Y(n2935_n), .Y(n2935) );
 INVXLTS U2289 ( .A(n2911), .A(n2911_n), .Y(n3562_n), .Y(n3562) );
 INVXLTS U2290 ( .A(n3370), .A(n3370_n), .Y(n3526_n), .Y(n3526) );
 AND2XLTS U2291 ( .A(n2890), .A(n2890_n), .B(n2909), .B(n2909_n), .Y(n3370_n), .Y(n3370) );
 NOR2XLTS U2292 ( .A(n3004), .A(n3004_n), .B(n2875), .B(n2875_n), .Y(n3003_n), .Y(n3003) );
 NOR2XLTS U2293 ( .A(n2866), .A(n2866_n), .B(n2883), .B(n2883_n), .Y(n3404_n), .Y(n3404) );
 NAND2X1TS U2294 ( .A(n3499), .A(n3499_n), .B(n3500), .B(n3500_n), .Y(n3131_n), .Y(n3131) );
 NOR2BX1TS U2295 ( .AN(n2906), .AN(n2906_n), .B(n2894), .B(n2894_n), .Y(n3500_n), .Y(n3500) );
 NOR2X1TS U2296 ( .A(n2902), .A(n2902_n), .B(n2900), .B(n2900_n), .Y(n3499_n), .Y(n3499) );
 NOR2BX1TS U2297 ( .AN(n2897), .AN(n2897_n), .B(n2913), .B(n2913_n), .Y(n3466_n), .Y(n3466) );
 NOR2BX1TS U2298 ( .AN(n2894), .AN(n2894_n), .B(n2905), .B(n2905_n), .Y(n3459_n), .Y(n3459) );
 NOR2BX1TS U2299 ( .AN(n2900), .AN(n2900_n), .B(n2902), .B(n2902_n), .Y(n3555_n), .Y(n3555) );
 NAND2X1TS U2300 ( .A(n2912), .A(n2912_n), .B(n2896), .B(n2896_n), .Y(n3556_n), .Y(n3556) );
 NOR2BX1TS U2301 ( .AN(n2903), .AN(n2903_n), .B(n2899), .B(n2899_n), .Y(n3460_n), .Y(n3460) );
 NAND2X1TS U2302 ( .A(n2890), .A(n2890_n), .B(n3570), .B(n3570_n), .Y(n3289_n), .Y(n3289) );
 NAND2X1TS U2303 ( .A(n3466), .A(n3466_n), .B(n2889), .B(n2889_n), .Y(n3465_n), .Y(n3465) );
 NAND2X1TS U2304 ( .A(n2961), .A(n2961_n), .B(n2962), .B(n2962_n), .Y(d[6]_n), .Y(d[6]) );
 NAND2X1TS U2305 ( .A(n2965), .A(n2965_n), .B(n2966), .B(n2966_n), .Y(n2964_n), .Y(n2964) );
 NAND2X1TS U2306 ( .A(n2969), .A(n2969_n), .B(n2970), .B(n2970_n), .Y(n2967_n), .Y(n2967) );
 NAND2X1TS U2307 ( .A(n2973), .A(n2973_n), .B(n2974), .B(n2974_n), .Y(n2972_n), .Y(n2972) );
 NAND2X1TS U2308 ( .A(n2870), .A(n2870_n), .B(n2738), .B(n2738_n), .Y(n2974_n), .Y(n2974) );
 NAND2X1TS U2309 ( .A(n2817), .A(n2817_n), .B(n2976), .B(n2976_n), .Y(n2973_n), .Y(n2973) );
 NAND2X1TS U2310 ( .A(n2980), .A(n2980_n), .B(n2981), .B(n2981_n), .Y(n2979_n), .Y(n2979) );
 NAND2BX1TS U2311 ( .AN(n2982), .AN(n2982_n), .B(n2810), .B(n2810_n), .Y(n2981_n), .Y(n2981) );
 NAND2X1TS U2312 ( .A(n2786), .A(n2786_n), .B(n2983), .B(n2983_n), .Y(n2980_n), .Y(n2980) );
 NAND2X1TS U2313 ( .A(n2780), .A(n2780_n), .B(n2758), .B(n2758_n), .Y(n2983_n), .Y(n2983) );
 NAND2X1TS U2314 ( .A(n2984), .A(n2984_n), .B(n2985), .B(n2985_n), .Y(n2978_n), .Y(n2978) );
 NAND2X1TS U2315 ( .A(n2859), .A(n2859_n), .B(n2987), .B(n2987_n), .Y(n2985_n), .Y(n2985) );
 NAND2X1TS U2316 ( .A(n2791), .A(n2791_n), .B(n2753), .B(n2753_n), .Y(n2987_n), .Y(n2987) );
 NAND2X1TS U2317 ( .A(n2844), .A(n2844_n), .B(n2989), .B(n2989_n), .Y(n2984_n), .Y(n2984) );
 NAND2X1TS U2318 ( .A(n2990), .A(n2990_n), .B(n2823), .B(n2823_n), .Y(n2989_n), .Y(n2989) );
 NAND2X1TS U2319 ( .A(n2992), .A(n2992_n), .B(n2993), .B(n2993_n), .Y(n2991_n), .Y(n2991) );
 NAND2X1TS U2320 ( .A(n2718), .A(n2718_n), .B(n2883), .B(n2883_n), .Y(n2993_n), .Y(n2993) );
 NAND2X1TS U2321 ( .A(n2994), .A(n2994_n), .B(n2769), .B(n2769_n), .Y(n2992_n), .Y(n2992) );
 NAND2X1TS U2322 ( .A(n3026), .A(n3026_n), .B(n3027), .B(n3027_n), .Y(d[5]_n), .Y(d[5]) );
 NAND2X1TS U2323 ( .A(n3030), .A(n3030_n), .B(n3031), .B(n3031_n), .Y(n3029_n), .Y(n3029) );
 NAND2X1TS U2324 ( .A(n3034), .A(n3034_n), .B(n3035), .B(n3035_n), .Y(n3033_n), .Y(n3033) );
 NAND2X1TS U2325 ( .A(n3041), .A(n3041_n), .B(n3042), .B(n3042_n), .Y(n3032_n), .Y(n3032) );
 NAND2X1TS U2326 ( .A(n2727), .A(n2727_n), .B(n3045), .B(n3045_n), .Y(n2976_n), .Y(n2976) );
 NAND2X1TS U2327 ( .A(n2908), .A(n2908_n), .B(n3046), .B(n3046_n), .Y(n3045_n), .Y(n3045) );
 NAND2X1TS U2328 ( .A(n3468), .A(n3468_n), .B(n3469), .B(n3469_n), .Y(n3467_n), .Y(n3467) );
 NAND2X1TS U2329 ( .A(n3472), .A(n3472_n), .B(n3473), .B(n3473_n), .Y(n3471_n), .Y(n3471) );
 NAND2X1TS U2330 ( .A(n2873), .A(n2873_n), .B(n2751), .B(n2751_n), .Y(n3473_n), .Y(n3473) );
 NAND2X1TS U2331 ( .A(n2852), .A(n2852_n), .B(n3424), .B(n3424_n), .Y(n3472_n), .Y(n3472) );
 NAND2X1TS U2332 ( .A(n3476), .A(n3476_n), .B(n3477), .B(n3477_n), .Y(n3475_n), .Y(n3475) );
 NAND2X1TS U2333 ( .A(n3051), .A(n3051_n), .B(n3156), .B(n3156_n), .Y(n3477_n), .Y(n3477) );
 NAND2X1TS U2334 ( .A(n2810), .A(n2810_n), .B(n3478), .B(n3478_n), .Y(n3476_n), .Y(n3476) );
 NAND2X1TS U2335 ( .A(n2834), .A(n2834_n), .B(n2768), .B(n2768_n), .Y(n3478_n), .Y(n3478) );
 NAND2X1TS U2336 ( .A(n3479), .A(n3479_n), .B(n3480), .B(n3480_n), .Y(n3474_n), .Y(n3474) );
 NAND2X1TS U2337 ( .A(n2870), .A(n2870_n), .B(n3481), .B(n3481_n), .Y(n3480_n), .Y(n3480) );
 NAND2X1TS U2338 ( .A(n2827), .A(n2827_n), .B(n3482), .B(n3482_n), .Y(n3481_n), .Y(n3481) );
 NAND2X1TS U2339 ( .A(n2906), .A(n2906_n), .B(n2709), .B(n2709_n), .Y(n3482_n), .Y(n3482) );
 NAND2X1TS U2340 ( .A(n3054), .A(n3054_n), .B(n3055), .B(n3055_n), .Y(n3052_n), .Y(n3052) );
 NAND2X1TS U2341 ( .A(n3060), .A(n3060_n), .B(n3061), .B(n3061_n), .Y(d[4]_n), .Y(d[4]) );
 NAND2X1TS U2342 ( .A(n3063), .A(n3063_n), .B(n3064), .B(n3064_n), .Y(n3062_n), .Y(n3062) );
 NOR2BX1TS U2343 ( .AN(n2951), .AN(n2951_n), .B(n3065), .B(n3065_n), .Y(n3064_n), .Y(n3064) );
 NAND2X1TS U2344 ( .A(n2959), .A(n2959_n), .B(n3066), .B(n3066_n), .Y(n3065_n), .Y(n3065) );
 NAND2X1TS U2345 ( .A(n3069), .A(n3069_n), .B(n3070), .B(n3070_n), .Y(n3068_n), .Y(n3068) );
 NAND2X1TS U2346 ( .A(n2845), .A(n2845_n), .B(n2859), .B(n2859_n), .Y(n3069_n), .Y(n3069) );
 NAND2X1TS U2347 ( .A(n3100), .A(n3100_n), .B(n3101), .B(n3101_n), .Y(n3099_n), .Y(n3099) );
 NAND2X1TS U2348 ( .A(n2747), .A(n2747_n), .B(n3102), .B(n3102_n), .Y(n3101_n), .Y(n3101) );
 NAND2X1TS U2349 ( .A(n2760), .A(n2760_n), .B(n2826), .B(n2826_n), .Y(n3102_n), .Y(n3102) );
 NAND2X1TS U2350 ( .A(n2754), .A(n2754_n), .B(n3103), .B(n3103_n), .Y(n3100_n), .Y(n3100) );
 NAND2X1TS U2351 ( .A(n3104), .A(n3104_n), .B(n2758), .B(n2758_n), .Y(n3103_n), .Y(n3103) );
 NAND2X1TS U2352 ( .A(n3105), .A(n3105_n), .B(n3106), .B(n3106_n), .Y(n3098_n), .Y(n3098) );
 NAND2X1TS U2353 ( .A(n3113), .A(n3113_n), .B(n3114), .B(n3114_n), .Y(n3112_n), .Y(n3112) );
 NAND2X1TS U2354 ( .A(n2726), .A(n2726_n), .B(n2786), .B(n2786_n), .Y(n3114_n), .Y(n3114) );
 NAND2X1TS U2355 ( .A(n2769), .A(n2769_n), .B(n3115), .B(n3115_n), .Y(n3113_n), .Y(n3113) );
 NAND2X1TS U2356 ( .A(n3117), .A(n3117_n), .B(n3118), .B(n3118_n), .Y(n3116_n), .Y(n3116) );
 NAND2X1TS U2357 ( .A(n3121), .A(n3121_n), .B(n3122), .B(n3122_n), .Y(n3120_n), .Y(n3120) );
 NAND2X1TS U2358 ( .A(n3128), .A(n3128_n), .B(n3129), .B(n3129_n), .Y(n3127_n), .Y(n3127) );
 NAND2X1TS U2359 ( .A(n2871), .A(n2871_n), .B(n3130), .B(n3130_n), .Y(n3129_n), .Y(n3129) );
 NAND2X1TS U2360 ( .A(n2821), .A(n2821_n), .B(n2724), .B(n2724_n), .Y(n3130_n), .Y(n3130) );
 NAND2X1TS U2361 ( .A(n2770), .A(n2770_n), .B(n3132), .B(n3132_n), .Y(n3128_n), .Y(n3128) );
 NAND2X1TS U2362 ( .A(n3139), .A(n3139_n), .B(n3140), .B(n3140_n), .Y(n3138_n), .Y(n3138) );
 NAND2X1TS U2363 ( .A(n2862), .A(n2862_n), .B(n2852), .B(n2852_n), .Y(n3140_n), .Y(n3140) );
 NAND2X1TS U2364 ( .A(n2748), .A(n2748_n), .B(n2785), .B(n2785_n), .Y(n3139_n), .Y(n3139) );
 NAND2X1TS U2365 ( .A(n3142), .A(n3142_n), .B(n3143), .B(n3143_n), .Y(n3137_n), .Y(n3137) );
 NAND2X1TS U2366 ( .A(n2755), .A(n2755_n), .B(n2779), .B(n2779_n), .Y(n3143_n), .Y(n3143) );
 NAND2X1TS U2367 ( .A(n2865), .A(n2865_n), .B(n2848), .B(n2848_n), .Y(n3142_n), .Y(n3142) );
 NAND2X1TS U2368 ( .A(n2914), .A(n2914_n), .B(n2915), .B(n2915_n), .Y(d[7]_n), .Y(d[7]) );
 NAND2X1TS U2369 ( .A(n2995), .A(n2995_n), .B(n2996), .B(n2996_n), .Y(n2917_n), .Y(n2917) );
 NAND2X1TS U2370 ( .A(n2999), .A(n2999_n), .B(n3000), .B(n3000_n), .Y(n2998_n), .Y(n2998) );
 NAND2X1TS U2371 ( .A(n3009), .A(n3009_n), .B(n3010), .B(n3010_n), .Y(n3008_n), .Y(n3008) );
 NAND2X1TS U2372 ( .A(n2725), .A(n2725_n), .B(n2713), .B(n2713_n), .Y(n3010_n), .Y(n3010) );
 NAND2X1TS U2373 ( .A(n3017), .A(n3017_n), .B(n3018), .B(n3018_n), .Y(n2997_n), .Y(n2997) );
 NAND2X1TS U2374 ( .A(n3021), .A(n3021_n), .B(n3022), .B(n3022_n), .Y(n3020_n), .Y(n3020) );
 NAND2X1TS U2375 ( .A(n2750), .A(n2750_n), .B(n2755), .B(n2755_n), .Y(n3022_n), .Y(n3022) );
 NAND2X1TS U2376 ( .A(n2918), .A(n2918_n), .B(n2919), .B(n2919_n), .Y(n2916_n), .Y(n2916) );
 NAND2X1TS U2377 ( .A(n2922), .A(n2922_n), .B(n2923), .B(n2923_n), .Y(n2921_n), .Y(n2921) );
 NAND2X1TS U2378 ( .A(n2729), .A(n2729_n), .B(n2817), .B(n2817_n), .Y(n2923_n), .Y(n2923) );
 NAND2X1TS U2379 ( .A(n2882), .A(n2882_n), .B(n2797), .B(n2797_n), .Y(n2922_n), .Y(n2922) );
 NAND2X1TS U2380 ( .A(n2926), .A(n2926_n), .B(n2927), .B(n2927_n), .Y(n2920_n), .Y(n2920) );
 NAND2X1TS U2381 ( .A(n2770), .A(n2770_n), .B(n2878), .B(n2878_n), .Y(n2927_n), .Y(n2927) );
 NAND2X1TS U2382 ( .A(n2811), .A(n2811_n), .B(n2702), .B(n2702_n), .Y(n2926_n), .Y(n2926) );
 NAND2X1TS U2383 ( .A(n2931), .A(n2931_n), .B(n2932), .B(n2932_n), .Y(n2930_n), .Y(n2930) );
 NAND2X1TS U2384 ( .A(n2863), .A(n2863_n), .B(n2934), .B(n2934_n), .Y(n2932_n), .Y(n2932) );
 NAND2X1TS U2385 ( .A(n2887), .A(n2887_n), .B(n2936), .B(n2936_n), .Y(n2931_n), .Y(n2931) );
 NAND2X1TS U2386 ( .A(n2937), .A(n2937_n), .B(n2938), .B(n2938_n), .Y(n2929_n), .Y(n2929) );
 NAND2X1TS U2387 ( .A(n2857), .A(n2857_n), .B(n2940), .B(n2940_n), .Y(n2938_n), .Y(n2938) );
 NAND2X1TS U2388 ( .A(n2941), .A(n2941_n), .B(n2791), .B(n2791_n), .Y(n2940_n), .Y(n2940) );
 NAND2X1TS U2389 ( .A(n2706), .A(n2706_n), .B(n2898), .B(n2898_n), .Y(n2947_n), .Y(n2947) );
 NAND2X1TS U2390 ( .A(n2950), .A(n2950_n), .B(n2951), .B(n2951_n), .Y(n2949_n), .Y(n2949) );
 NAND2X1TS U2391 ( .A(n3083), .A(n3083_n), .B(n3084), .B(n3084_n), .Y(n3082_n), .Y(n3082) );
 NAND2X1TS U2392 ( .A(n2816), .A(n2816_n), .B(n2778), .B(n2778_n), .Y(n3084_n), .Y(n3084) );
 NAND2X1TS U2393 ( .A(n3090), .A(n3090_n), .B(n3091), .B(n3091_n), .Y(n3081_n), .Y(n3081) );
 NAND2X1TS U2394 ( .A(n2845), .A(n2845_n), .B(n3092), .B(n3092_n), .Y(n3091_n), .Y(n3091) );
 NAND2X1TS U2395 ( .A(n2712), .A(n2712_n), .B(n2720), .B(n2720_n), .Y(n3092_n), .Y(n3092) );
 NAND2X1TS U2396 ( .A(n3144), .A(n3144_n), .B(n3145), .B(n3145_n), .Y(n2953_n), .Y(n2953) );
 NAND2X1TS U2397 ( .A(n3148), .A(n3148_n), .B(n3149), .B(n3149_n), .Y(n3147_n), .Y(n3147) );
 NAND2X1TS U2398 ( .A(n2875), .A(n2875_n), .B(n3150), .B(n3150_n), .Y(n3149_n), .Y(n3149) );
 NAND2X1TS U2399 ( .A(n2811), .A(n2811_n), .B(n2745), .B(n2745_n), .Y(n3148_n), .Y(n3148) );
 NAND2X1TS U2400 ( .A(n3154), .A(n3154_n), .B(n3155), .B(n3155_n), .Y(n3153_n), .Y(n3153) );
 NAND2X1TS U2401 ( .A(n2784), .A(n2784_n), .B(n3156), .B(n3156_n), .Y(n3155_n), .Y(n3155) );
 NAND2X1TS U2402 ( .A(n2954), .A(n2954_n), .B(n2781), .B(n2781_n), .Y(n3156_n), .Y(n3156) );
 NAND2X1TS U2403 ( .A(n2787), .A(n2787_n), .B(n3157), .B(n3157_n), .Y(n3154_n), .Y(n3154) );
 NAND2X1TS U2404 ( .A(n3158), .A(n3158_n), .B(n2727), .B(n2727_n), .Y(n3157_n), .Y(n3157) );
 NAND2X1TS U2405 ( .A(n3159), .A(n3159_n), .B(n3160), .B(n3160_n), .Y(n3152_n), .Y(n3152) );
 NAND2X1TS U2406 ( .A(n2855), .A(n2855_n), .B(n3162), .B(n3162_n), .Y(n3160_n), .Y(n3160) );
 NAND2X1TS U2407 ( .A(n2982), .A(n2982_n), .B(n2721), .B(n2721_n), .Y(n3162_n), .Y(n3162) );
 NAND2X1TS U2408 ( .A(n2879), .A(n2879_n), .B(n3163), .B(n3163_n), .Y(n3159_n), .Y(n3159) );
 NAND2X1TS U2409 ( .A(n2796), .A(n2796_n), .B(n2789), .B(n2789_n), .Y(n3163_n), .Y(n3163) );
 NAND2X1TS U2410 ( .A(n2955), .A(n2955_n), .B(n2956), .B(n2956_n), .Y(n2948_n), .Y(n2948) );
 NAND2X1TS U2411 ( .A(n2959), .A(n2959_n), .B(n2960), .B(n2960_n), .Y(n2958_n), .Y(n2958) );
 NAND2X1TS U2412 ( .A(n3073), .A(n3073_n), .B(n3074), .B(n3074_n), .Y(n3072_n), .Y(n3072) );
 NAND2X1TS U2413 ( .A(n2885), .A(n2885_n), .B(n2849), .B(n2849_n), .Y(n3074_n), .Y(n3074) );
 NAND2X1TS U2414 ( .A(n2798), .A(n2798_n), .B(n2725), .B(n2725_n), .Y(n3073_n), .Y(n3073) );
 NAND2X1TS U2415 ( .A(n3075), .A(n3075_n), .B(n3076), .B(n3076_n), .Y(n3071_n), .Y(n3071) );
 NAND2X1TS U2416 ( .A(n2865), .A(n2865_n), .B(n2842), .B(n2842_n), .Y(n3076_n), .Y(n3076) );
 NAND2X1TS U2417 ( .A(n3510), .A(n3510_n), .B(n3511), .B(n3511_n), .Y(n3509_n), .Y(n3509) );
 NAND2X1TS U2418 ( .A(n3514), .A(n3514_n), .B(n3515), .B(n3515_n), .Y(n3513_n), .Y(n3513) );
 NAND2X1TS U2419 ( .A(n2855), .A(n2855_n), .B(n3257), .B(n3257_n), .Y(n3515_n), .Y(n3515) );
 NAND2X1TS U2420 ( .A(n3521), .A(n3521_n), .B(n3522), .B(n3522_n), .Y(n3520_n), .Y(n3520) );
 NAND2X1TS U2421 ( .A(n2816), .A(n2816_n), .B(n2874), .B(n2874_n), .Y(n3522_n), .Y(n3522) );
 NAND2X1TS U2422 ( .A(n2869), .A(n2869_n), .B(n3458), .B(n3458_n), .Y(n3521_n), .Y(n3521) );
 NAND2X1TS U2423 ( .A(n3528), .A(n3528_n), .B(n3529), .B(n3529_n), .Y(n3057_n), .Y(n3057) );
 NAND2X1TS U2424 ( .A(n3535), .A(n3535_n), .B(n3342), .B(n3342_n), .Y(n3534_n), .Y(n3534) );
 NAND2X1TS U2425 ( .A(n2766), .A(n2766_n), .B(n2822), .B(n2822_n), .Y(n3136_n), .Y(n3136) );
 NAND2X1TS U2426 ( .A(n3169), .A(n3169_n), .B(n2788), .B(n2788_n), .Y(n3168_n), .Y(n3168) );
 NAND2X1TS U2427 ( .A(n2753), .A(n2753_n), .B(n2736), .B(n2736_n), .Y(n3170_n), .Y(n3170) );
 NAND2X1TS U2428 ( .A(n2717), .A(n2717_n), .B(n2887), .B(n2887_n), .Y(n3070_n), .Y(n3070) );
 NAND2X1TS U2429 ( .A(n3173), .A(n3173_n), .B(n3174), .B(n3174_n), .Y(n3028_n), .Y(n3028) );
 NAND2X1TS U2430 ( .A(n3430), .A(n3430_n), .B(n3431), .B(n3431_n), .Y(n3176_n), .Y(n3176) );
 NAND2X1TS U2431 ( .A(n2747), .A(n2747_n), .B(n2713), .B(n2713_n), .Y(n3431_n), .Y(n3431) );
 NAND2X1TS U2432 ( .A(n3434), .A(n3434_n), .B(n3435), .B(n3435_n), .Y(n3433_n), .Y(n3433) );
 NAND2X1TS U2433 ( .A(n2863), .A(n2863_n), .B(n2787), .B(n2787_n), .Y(n3435_n), .Y(n3435) );
 NAND2X1TS U2434 ( .A(n2797), .A(n2797_n), .B(n2860), .B(n2860_n), .Y(n3434_n), .Y(n3434) );
 NAND2X1TS U2435 ( .A(n3436), .A(n3436_n), .B(n3437), .B(n3437_n), .Y(n3432_n), .Y(n3432) );
 NAND2X1TS U2436 ( .A(n2924), .A(n2924_n), .B(n2866), .B(n2866_n), .Y(n3437_n), .Y(n3437) );
 NAND2X1TS U2437 ( .A(n2754), .A(n2754_n), .B(n2882), .B(n2882_n), .Y(n3436_n), .Y(n3436) );
 NAND2X1TS U2438 ( .A(n3177), .A(n3177_n), .B(n3178), .B(n3178_n), .Y(n3175_n), .Y(n3175) );
 NAND2X1TS U2439 ( .A(n3181), .A(n3181_n), .B(n3182), .B(n3182_n), .Y(n3180_n), .Y(n3180) );
 NAND2X1TS U2440 ( .A(n2885), .A(n2885_n), .B(n3183), .B(n3183_n), .Y(n3182_n), .Y(n3182) );
 NAND2X1TS U2441 ( .A(n3191), .A(n3191_n), .B(n3192), .B(n3192_n), .Y(n3190_n), .Y(n3190) );
 NAND2X1TS U2442 ( .A(n2939), .A(n2939_n), .B(n3193), .B(n3193_n), .Y(n3192_n), .Y(n3192) );
 NAND2X1TS U2443 ( .A(n2795), .A(n2795_n), .B(n2803), .B(n2803_n), .Y(n3193_n), .Y(n3193) );
 NAND2X1TS U2444 ( .A(n2867), .A(n2867_n), .B(n3194), .B(n3194_n), .Y(n3191_n), .Y(n3191) );
 NAND2X1TS U2445 ( .A(n2820), .A(n2820_n), .B(n2775), .B(n2775_n), .Y(n3194_n), .Y(n3194) );
 NAND2X1TS U2446 ( .A(n3198), .A(n3198_n), .B(n3199), .B(n3199_n), .Y(n3197_n), .Y(n3197) );
 NAND2X1TS U2447 ( .A(n2849), .A(n2849_n), .B(n2870), .B(n2870_n), .Y(n3199_n), .Y(n3199) );
 NAND2X1TS U2448 ( .A(n3204), .A(n3204_n), .B(n3205), .B(n3205_n), .Y(n3179_n), .Y(n3179) );
 NAND2X1TS U2449 ( .A(n3209), .A(n3209_n), .B(n3210), .B(n3210_n), .Y(n3196_n), .Y(n3196) );
 NAND2X1TS U2450 ( .A(n2800), .A(n2800_n), .B(n2743), .B(n2743_n), .Y(n3166_n), .Y(n3166) );
 NAND2X1TS U2451 ( .A(n3216), .A(n3216_n), .B(n3217), .B(n3217_n), .Y(n3215_n), .Y(n3215) );
 NAND2BX1TS U2452 ( .AN(n2941), .AN(n2941_n), .B(n2860), .B(n2860_n), .Y(n3217_n), .Y(n3217) );
 NAND2X1TS U2453 ( .A(n2854), .A(n2854_n), .B(n3115), .B(n3115_n), .Y(n3216_n), .Y(n3216) );
 NAND2X1TS U2454 ( .A(n3487), .A(n3487_n), .B(n3488), .B(n3488_n), .Y(n3203_n), .Y(n3203) );
 NAND2X1TS U2455 ( .A(n3490), .A(n3490_n), .B(n3491), .B(n3491_n), .Y(n3489_n), .Y(n3489) );
 NAND2X1TS U2456 ( .A(n2817), .A(n2817_n), .B(n2886), .B(n2886_n), .Y(n3491_n), .Y(n3491) );
 NAND2X1TS U2457 ( .A(n3496), .A(n3496_n), .B(n3497), .B(n3497_n), .Y(n3495_n), .Y(n3495) );
 NAND2X1TS U2458 ( .A(n3004), .A(n3004_n), .B(n3150), .B(n3150_n), .Y(n3497_n), .Y(n3497) );
 NAND2X1TS U2459 ( .A(n3498), .A(n3498_n), .B(n2804), .B(n2804_n), .Y(n3150_n), .Y(n3150) );
 NAND2BX1TS U2460 ( .AN(n3384), .AN(n3384_n), .B(n2852), .B(n2852_n), .Y(n3496_n), .Y(n3496) );
 NAND2X1TS U2461 ( .A(n3501), .A(n3501_n), .B(n3502), .B(n3502_n), .Y(n3494_n), .Y(n3494) );
 NAND2X1TS U2462 ( .A(n2730), .A(n2730_n), .B(n3503), .B(n3503_n), .Y(n3502_n), .Y(n3502) );
 NAND2X1TS U2463 ( .A(n3047), .A(n3047_n), .B(n2771), .B(n2771_n), .Y(n3503_n), .Y(n3503) );
 NAND2X1TS U2464 ( .A(n2885), .A(n2885_n), .B(n2783), .B(n2783_n), .Y(n3220_n), .Y(n3220) );
 NAND2X1TS U2465 ( .A(n2755), .A(n2755_n), .B(n2879), .B(n2879_n), .Y(n3219_n), .Y(n3219) );
 NAND2X1TS U2466 ( .A(n3109), .A(n3109_n), .B(n3222), .B(n3222_n), .Y(n3221_n), .Y(n3221) );
 NAND2X1TS U2467 ( .A(n2790), .A(n2790_n), .B(n2774), .B(n2774_n), .Y(n2934_n), .Y(n2934) );
 NAND2X1TS U2468 ( .A(n3228), .A(n3228_n), .B(n3229), .B(n3229_n), .Y(n3227_n), .Y(n3227) );
 NAND2X1TS U2469 ( .A(n3006), .A(n3006_n), .B(n2936), .B(n2936_n), .Y(n3229_n), .Y(n3229) );
 NAND2X1TS U2470 ( .A(n2988), .A(n2988_n), .B(n2731), .B(n2731_n), .Y(n2936_n), .Y(n2936) );
 NAND2X1TS U2471 ( .A(n3232), .A(n3232_n), .B(n3233), .B(n3233_n), .Y(n3231_n), .Y(n3231) );
 NAND2BX1TS U2472 ( .AN(n3088), .AN(n3088_n), .B(n2765), .B(n2765_n), .Y(n3233_n), .Y(n3233) );
 NAND2X1TS U2473 ( .A(n2844), .A(n2844_n), .B(n3234), .B(n3234_n), .Y(n3232_n), .Y(n3232) );
 NAND2X1TS U2474 ( .A(n2782), .A(n2782_n), .B(n2716), .B(n2716_n), .Y(n3234_n), .Y(n3234) );
 NAND2X1TS U2475 ( .A(n3236), .A(n3236_n), .B(n3237), .B(n3237_n), .Y(n3226_n), .Y(n3226) );
 NAND2X1TS U2476 ( .A(n3240), .A(n3240_n), .B(n3241), .B(n3241_n), .Y(n3239_n), .Y(n3239) );
 NAND2X1TS U2477 ( .A(n2729), .A(n2729_n), .B(n2784), .B(n2784_n), .Y(n3241_n), .Y(n3241) );
 NAND2X1TS U2478 ( .A(n3242), .A(n3242_n), .B(n3243), .B(n3243_n), .Y(n3238_n), .Y(n3238) );
 NAND2X1TS U2479 ( .A(n2888), .A(n2888_n), .B(n2810), .B(n2810_n), .Y(n3243_n), .Y(n3243) );
 NAND2X1TS U2480 ( .A(n3004), .A(n3004_n), .B(n2770), .B(n2770_n), .Y(n3245_n), .Y(n3245) );
 NAND2X1TS U2481 ( .A(n3442), .A(n3442_n), .B(n3443), .B(n3443_n), .Y(n3441_n), .Y(n3441) );
 NAND2X1TS U2482 ( .A(n2883), .A(n2883_n), .B(n2737), .B(n2737_n), .Y(n3443_n), .Y(n3443) );
 NAND2X1TS U2483 ( .A(n2770), .A(n2770_n), .B(n3330), .B(n3330_n), .Y(n3442_n), .Y(n3442) );
 NAND2X1TS U2484 ( .A(n3444), .A(n3444_n), .B(n3445), .B(n3445_n), .Y(n3440_n), .Y(n3440) );
 NAND2X1TS U2485 ( .A(n3446), .A(n3446_n), .B(n2764), .B(n2764_n), .Y(n3445_n), .Y(n3445) );
 NAND2X1TS U2486 ( .A(n2862), .A(n2862_n), .B(n3447), .B(n3447_n), .Y(n3444_n), .Y(n3444) );
 NAND2X1TS U2487 ( .A(n2819), .A(n2819_n), .B(n2840), .B(n2840_n), .Y(n3447_n), .Y(n3447) );
 NAND2X1TS U2488 ( .A(n3448), .A(n3448_n), .B(n3449), .B(n3449_n), .Y(n3438_n), .Y(n3438) );
 NAND2X1TS U2489 ( .A(n3454), .A(n3454_n), .B(n3455), .B(n3455_n), .Y(n3453_n), .Y(n3453) );
 NAND2X1TS U2490 ( .A(n2887), .A(n2887_n), .B(n2785), .B(n2785_n), .Y(n3455_n), .Y(n3455) );
 NAND2X1TS U2491 ( .A(n3249), .A(n3249_n), .B(n3250), .B(n3250_n), .Y(n3165_n), .Y(n3165) );
 NAND2X1TS U2492 ( .A(n3253), .A(n3253_n), .B(n3254), .B(n3254_n), .Y(n3252_n), .Y(n3252) );
 NAND2X1TS U2493 ( .A(n2750), .A(n2750_n), .B(n2809), .B(n2809_n), .Y(n3254_n), .Y(n3254) );
 NAND2X1TS U2494 ( .A(n2875), .A(n2875_n), .B(n2714), .B(n2714_n), .Y(n3253_n), .Y(n3253) );
 NAND2X1TS U2495 ( .A(n3255), .A(n3255_n), .B(n3256), .B(n3256_n), .Y(n3251_n), .Y(n3251) );
 NAND2X1TS U2496 ( .A(n2754), .A(n2754_n), .B(n3257), .B(n3257_n), .Y(n3256_n), .Y(n3256) );
 NAND2X1TS U2497 ( .A(n2860), .A(n2860_n), .B(n3258), .B(n3258_n), .Y(n3255_n), .Y(n3255) );
 NAND2X1TS U2498 ( .A(n3261), .A(n3261_n), .B(n3262), .B(n3262_n), .Y(n3260_n), .Y(n3260) );
 NAND2X1TS U2499 ( .A(n2763), .A(n2763_n), .B(n3263), .B(n3263_n), .Y(n3262_n), .Y(n3262) );
 NAND2X1TS U2500 ( .A(n3040), .A(n3040_n), .B(n2782), .B(n2782_n), .Y(n3263_n), .Y(n3263) );
 NAND2X1TS U2501 ( .A(n3006), .A(n3006_n), .B(n3264), .B(n3264_n), .Y(n3261_n), .Y(n3261) );
 NAND2X1TS U2502 ( .A(n2792), .A(n2792_n), .B(n2776), .B(n2776_n), .Y(n3264_n), .Y(n3264) );
 NAND2X1TS U2503 ( .A(n3265), .A(n3265_n), .B(n3266), .B(n3266_n), .Y(n3259_n), .Y(n3259) );
 NAND2X1TS U2504 ( .A(n2751), .A(n2751_n), .B(n3267), .B(n3267_n), .Y(n3266_n), .Y(n3266) );
 NAND2X1TS U2505 ( .A(n2711), .A(n2711_n), .B(n2721), .B(n2721_n), .Y(n3267_n), .Y(n3267) );
 NAND2X1TS U2506 ( .A(n2886), .A(n2886_n), .B(n3268), .B(n3268_n), .Y(n3265_n), .Y(n3265) );
 NAND2X1TS U2507 ( .A(n2805), .A(n2805_n), .B(n2828), .B(n2828_n), .Y(n3268_n), .Y(n3268) );
 NAND2X1TS U2508 ( .A(n3538), .A(n3538_n), .B(n3539), .B(n3539_n), .Y(n3247_n), .Y(n3247) );
 NAND2X1TS U2509 ( .A(n3541), .A(n3541_n), .B(n3542), .B(n3542_n), .Y(n3540_n), .Y(n3540) );
 NAND2X1TS U2510 ( .A(n2756), .A(n2756_n), .B(n3543), .B(n3543_n), .Y(n3542_n), .Y(n3542) );
 NAND2X1TS U2511 ( .A(n3544), .A(n3544_n), .B(n2833), .B(n2833_n), .Y(n3543_n), .Y(n3543) );
 NAND2X1TS U2512 ( .A(n3547), .A(n3547_n), .B(n3548), .B(n3548_n), .Y(n3546_n), .Y(n3546) );
 NAND2X1TS U2513 ( .A(n2783), .A(n2783_n), .B(n3549), .B(n3549_n), .Y(n3548_n), .Y(n3548) );
 NAND2X1TS U2514 ( .A(n2739), .A(n2739_n), .B(n2767), .B(n2767_n), .Y(n3549_n), .Y(n3549) );
 NAND2X1TS U2515 ( .A(n2846), .A(n2846_n), .B(n3550), .B(n3550_n), .Y(n3547_n), .Y(n3547) );
 NAND2X1TS U2516 ( .A(n3040), .A(n3040_n), .B(n2733), .B(n2733_n), .Y(n3550_n), .Y(n3550) );
 NAND2X1TS U2517 ( .A(n2839), .A(n2839_n), .B(n2759), .B(n2759_n), .Y(n3134_n), .Y(n3134) );
 NAND2X1TS U2518 ( .A(n3551), .A(n3551_n), .B(n3552), .B(n3552_n), .Y(n3545_n), .Y(n3545) );
 NAND2X1TS U2519 ( .A(n2925), .A(n2925_n), .B(n3553), .B(n3553_n), .Y(n3552_n), .Y(n3552) );
 NAND2X1TS U2520 ( .A(n3169), .A(n3169_n), .B(n2775), .B(n2775_n), .Y(n3553_n), .Y(n3553) );
 NAND2X1TS U2521 ( .A(n2866), .A(n2866_n), .B(n3554), .B(n3554_n), .Y(n3551_n), .Y(n3551) );
 NAND2X1TS U2522 ( .A(n2732), .A(n2732_n), .B(n2827), .B(n2827_n), .Y(n3554_n), .Y(n3554) );
 NAND2X1TS U2523 ( .A(n3557), .A(n3557_n), .B(n3558), .B(n3558_n), .Y(n3059_n), .Y(n3059) );
 NAND2X1TS U2524 ( .A(n3097), .A(n3097_n), .B(n3559), .B(n3559_n), .Y(n3558_n), .Y(n3558) );
 NAND2X1TS U2525 ( .A(n3544), .A(n3544_n), .B(n2839), .B(n2839_n), .Y(n3559_n), .Y(n3559) );
 NAND2X1TS U2526 ( .A(n3566), .A(n3566_n), .B(n3567), .B(n3567_n), .Y(n3565_n), .Y(n3565) );
 NAND2X1TS U2527 ( .A(n2756), .A(n2756_n), .B(n3464), .B(n3464_n), .Y(n3567_n), .Y(n3567) );
 NAND2X1TS U2528 ( .A(n3015), .A(n3015_n), .B(n2766), .B(n2766_n), .Y(n3464_n), .Y(n3464) );
 NAND2X1TS U2529 ( .A(n3023), .A(n3023_n), .B(n3571), .B(n3571_n), .Y(n3566_n), .Y(n3566) );
 NAND2X1TS U2530 ( .A(n2803), .A(n2803_n), .B(n2752), .B(n2752_n), .Y(n3571_n), .Y(n3571) );
 NAND2X1TS U2531 ( .A(n2774), .A(n2774_n), .B(n2735), .B(n2735_n), .Y(n3574_n), .Y(n3574) );
 NAND2X1TS U2532 ( .A(n3576), .A(n3576_n), .B(n3577), .B(n3577_n), .Y(n3575_n), .Y(n3575) );
 NAND2X1TS U2533 ( .A(n2888), .A(n2888_n), .B(n2797), .B(n2797_n), .Y(n3577_n), .Y(n3577) );
 NAND2X1TS U2534 ( .A(n2858), .A(n2858_n), .B(n3579), .B(n3579_n), .Y(n3576_n), .Y(n3576) );
 NAND2X1TS U2535 ( .A(n2761), .A(n2761_n), .B(n2814), .B(n2814_n), .Y(n3579_n), .Y(n3579) );
 NAND2X1TS U2536 ( .A(n3580), .A(n3580_n), .B(n3581), .B(n3581_n), .Y(n3058_n), .Y(n3058) );
 NAND2X1TS U2537 ( .A(n3060), .A(n3060_n), .B(n3269), .B(n3269_n), .Y(d[1]_n), .Y(d[1]) );
 NAND2X1TS U2538 ( .A(n3272), .A(n3272_n), .B(n3273), .B(n3273_n), .Y(n3271_n), .Y(n3271) );
 NAND2X1TS U2539 ( .A(n3274), .A(n3274_n), .B(n3275), .B(n3275_n), .Y(n2968_n), .Y(n2968) );
 NAND2X1TS U2540 ( .A(n3278), .A(n3278_n), .B(n3279), .B(n3279_n), .Y(n3277_n), .Y(n3277) );
 NAND2X1TS U2541 ( .A(n2867), .A(n2867_n), .B(n2798), .B(n2798_n), .Y(n3279_n), .Y(n3279) );
 NAND2X1TS U2542 ( .A(n2846), .A(n2846_n), .B(n2877), .B(n2877_n), .Y(n3278_n), .Y(n3278) );
 NAND2X1TS U2543 ( .A(n3280), .A(n3280_n), .B(n3281), .B(n3281_n), .Y(n3276_n), .Y(n3276) );
 NAND2X1TS U2544 ( .A(n2764), .A(n2764_n), .B(n2881), .B(n2881_n), .Y(n3281_n), .Y(n3281) );
 NAND2X1TS U2545 ( .A(n3285), .A(n3285_n), .B(n3286), .B(n3286_n), .Y(n3284_n), .Y(n3284) );
 NAND2X1TS U2546 ( .A(n2848), .A(n2848_n), .B(n3287), .B(n3287_n), .Y(n3286_n), .Y(n3286) );
 NAND2X1TS U2547 ( .A(n3104), .A(n3104_n), .B(n2739), .B(n2739_n), .Y(n3287_n), .Y(n3287) );
 NAND2X1TS U2548 ( .A(n3161), .A(n3161_n), .B(n3132), .B(n3132_n), .Y(n3285_n), .Y(n3285) );
 NAND2X1TS U2549 ( .A(n3290), .A(n3290_n), .B(n3291), .B(n3291_n), .Y(n3283_n), .Y(n3283) );
 NAND2X1TS U2550 ( .A(n2841), .A(n2841_n), .B(n3292), .B(n3292_n), .Y(n3291_n), .Y(n3291) );
 NAND2X1TS U2551 ( .A(n2837), .A(n2837_n), .B(n2823), .B(n2823_n), .Y(n3292_n), .Y(n3292) );
 NAND2X1TS U2552 ( .A(n3296), .A(n3296_n), .B(n3297), .B(n3297_n), .Y(n2957_n), .Y(n2957) );
 NAND2X1TS U2553 ( .A(n3302), .A(n3302_n), .B(n3303), .B(n3303_n), .Y(n3301_n), .Y(n3301) );
 NAND2X1TS U2554 ( .A(n3304), .A(n3304_n), .B(n2878), .B(n2878_n), .Y(n3303_n), .Y(n3303) );
 NAND2X1TS U2555 ( .A(n2765), .A(n2765_n), .B(n2986), .B(n2986_n), .Y(n3302_n), .Y(n3302) );
 NAND2X1TS U2556 ( .A(n3307), .A(n3307_n), .B(n3308), .B(n3308_n), .Y(n3306_n), .Y(n3306) );
 NAND2X1TS U2557 ( .A(n3313), .A(n3313_n), .B(n3314), .B(n3314_n), .Y(n3305_n), .Y(n3305) );
 NAND2X1TS U2558 ( .A(n2781), .A(n2781_n), .B(n2728), .B(n2728_n), .Y(n3257_n), .Y(n3257) );
 NAND2X1TS U2559 ( .A(n2960), .A(n2960_n), .B(n3323), .B(n3323_n), .Y(n3322_n), .Y(n3322) );
 NAND2X1TS U2560 ( .A(n3328), .A(n3328_n), .B(n3329), .B(n3329_n), .Y(n3327_n), .Y(n3327) );
 NAND2X1TS U2561 ( .A(n2701), .A(n2701_n), .B(n2737), .B(n2737_n), .Y(n3329_n), .Y(n3329) );
 NAND2X1TS U2562 ( .A(n2854), .A(n2854_n), .B(n3330), .B(n3330_n), .Y(n3328_n), .Y(n3328) );
 NAND2X1TS U2563 ( .A(n3331), .A(n3331_n), .B(n3332), .B(n3332_n), .Y(n3326_n), .Y(n3326) );
 NAND2X1TS U2564 ( .A(n2858), .A(n2858_n), .B(n3333), .B(n3333_n), .Y(n3332_n), .Y(n3332) );
 NAND2X1TS U2565 ( .A(n2977), .A(n2977_n), .B(n2830), .B(n2830_n), .Y(n3333_n), .Y(n3333) );
 NAND2X1TS U2566 ( .A(n3338), .A(n3338_n), .B(n3339), .B(n3339_n), .Y(n3019_n), .Y(n3019) );
 NAND2X1TS U2567 ( .A(n3240), .A(n3240_n), .B(n3342), .B(n3342_n), .Y(n3341_n), .Y(n3341) );
 NAND2X1TS U2568 ( .A(n2886), .A(n2886_n), .B(n2769), .B(n2769_n), .Y(n3342_n), .Y(n3342) );
 NAND2X1TS U2569 ( .A(n3023), .A(n3023_n), .B(n2786), .B(n2786_n), .Y(n3240_n), .Y(n3240) );
 NAND2X1TS U2570 ( .A(n3343), .A(n3343_n), .B(n3344), .B(n3344_n), .Y(n3340_n), .Y(n3340) );
 NAND2X1TS U2571 ( .A(n3097), .A(n3097_n), .B(n3330), .B(n3330_n), .Y(n3344_n), .Y(n3344) );
 NAND2X1TS U2572 ( .A(n2704), .A(n2704_n), .B(n2742), .B(n2742_n), .Y(n3330_n), .Y(n3330) );
 NAND2X1TS U2573 ( .A(n2857), .A(n2857_n), .B(n2763), .B(n2763_n), .Y(n3343_n), .Y(n3343) );
 NAND2X1TS U2574 ( .A(n3347), .A(n3347_n), .B(n3348), .B(n3348_n), .Y(n3346_n), .Y(n3346) );
 NAND2X1TS U2575 ( .A(n2809), .A(n2809_n), .B(n3349), .B(n3349_n), .Y(n3348_n), .Y(n3348) );
 NAND2X1TS U2576 ( .A(n3350), .A(n3350_n), .B(n2781), .B(n2781_n), .Y(n3349_n), .Y(n3349) );
 NAND2X1TS U2577 ( .A(n2877), .A(n2877_n), .B(n3351), .B(n3351_n), .Y(n3347_n), .Y(n3347) );
 NAND2X1TS U2578 ( .A(n3169), .A(n3169_n), .B(n2802), .B(n2802_n), .Y(n3351_n), .Y(n3351) );
 NAND2X1TS U2579 ( .A(n3352), .A(n3352_n), .B(n3353), .B(n3353_n), .Y(n3345_n), .Y(n3345) );
 NAND2X1TS U2580 ( .A(n2924), .A(n2924_n), .B(n3354), .B(n3354_n), .Y(n3353_n), .Y(n3353) );
 NAND2X1TS U2581 ( .A(n2838), .A(n2838_n), .B(n2767), .B(n2767_n), .Y(n3354_n), .Y(n3354) );
 NAND2X1TS U2582 ( .A(n2744), .A(n2744_n), .B(n3355), .B(n3355_n), .Y(n3352_n), .Y(n3352) );
 NAND2X1TS U2583 ( .A(n3295), .A(n3295_n), .B(n2831), .B(n2831_n), .Y(n3355_n), .Y(n3355) );
 NAND2X1TS U2584 ( .A(n2707), .A(n2707_n), .B(n3460), .B(n3460_n), .Y(n3013_n), .Y(n3013) );
 NAND2X1TS U2585 ( .A(n2820), .A(n2820_n), .B(n2792), .B(n2792_n), .Y(n3356_n), .Y(n3356) );
 NAND2X1TS U2586 ( .A(n3359), .A(n3359_n), .B(n3360), .B(n3360_n), .Y(n3358_n), .Y(n3358) );
 NAND2X1TS U2587 ( .A(n2798), .A(n2798_n), .B(n3361), .B(n3361_n), .Y(n3360_n), .Y(n3360) );
 NAND2X1TS U2588 ( .A(n2800), .A(n2800_n), .B(n2757), .B(n2757_n), .Y(n3361_n), .Y(n3361) );
 NAND2X1TS U2589 ( .A(n2911), .A(n2911_n), .B(n2908), .B(n2908_n), .Y(n3573_n), .Y(n3573) );
 NAND2X1TS U2590 ( .A(n2726), .A(n2726_n), .B(n3362), .B(n3362_n), .Y(n3359_n), .Y(n3359) );
 NAND2X1TS U2591 ( .A(n2829), .A(n2829_n), .B(n2735), .B(n2735_n), .Y(n3362_n), .Y(n3362) );
 NAND2X1TS U2592 ( .A(n3366), .A(n3366_n), .B(n3367), .B(n3367_n), .Y(n3365_n), .Y(n3365) );
 NAND2X1TS U2593 ( .A(n2844), .A(n2844_n), .B(n2865), .B(n2865_n), .Y(n3367_n), .Y(n3367) );
 NAND2X1TS U2594 ( .A(n3370), .A(n3370_n), .B(n2897), .B(n2897_n), .Y(n3167_n), .Y(n3167) );
 NAND2X1TS U2595 ( .A(n3373), .A(n3373_n), .B(n3374), .B(n3374_n), .Y(n3372_n), .Y(n3372) );
 NAND2X1TS U2596 ( .A(n3499), .A(n3499_n), .B(n2706), .B(n2706_n), .Y(n2988_n), .Y(n2988) );
 NAND2X1TS U2597 ( .A(n3379), .A(n3379_n), .B(n3244), .B(n3244_n), .Y(n3378_n), .Y(n3378) );
 NAND2X1TS U2598 ( .A(n2869), .A(n2869_n), .B(n2851), .B(n2851_n), .Y(n3244_n), .Y(n3244) );
 NAND2X1TS U2599 ( .A(n2881), .A(n2881_n), .B(n2848), .B(n2848_n), .Y(n3379_n), .Y(n3379) );
 NAND2X1TS U2600 ( .A(n3459), .A(n3459_n), .B(n2709), .B(n2709_n), .Y(n3125_n), .Y(n3125) );
 NAND2X1TS U2601 ( .A(n3380), .A(n3380_n), .B(n3381), .B(n3381_n), .Y(n3371_n), .Y(n3371) );
 NAND2X1TS U2602 ( .A(n3387), .A(n3387_n), .B(n3388), .B(n3388_n), .Y(n3386_n), .Y(n3386) );
 NAND2X1TS U2603 ( .A(n2866), .A(n2866_n), .B(n3389), .B(n3389_n), .Y(n3388_n), .Y(n3388) );
 NAND2X1TS U2604 ( .A(n2794), .A(n2794_n), .B(n2829), .B(n2829_n), .Y(n3389_n), .Y(n3389) );
 NAND2X1TS U2605 ( .A(n3459), .A(n3459_n), .B(n3428), .B(n3428_n), .Y(n3089_n), .Y(n3089) );
 NAND2X1TS U2606 ( .A(n2874), .A(n2874_n), .B(n3258), .B(n3258_n), .Y(n3387_n), .Y(n3387) );
 NAND2X1TS U2607 ( .A(n2795), .A(n2795_n), .B(n2723), .B(n2723_n), .Y(n3258_n), .Y(n3258) );
 NAND2X1TS U2608 ( .A(n2740), .A(n2740_n), .B(n2838), .B(n2838_n), .Y(n3115_n), .Y(n3115) );
 NAND2X1TS U2609 ( .A(n2730), .A(n2730_n), .B(n2845), .B(n2845_n), .Y(n3391_n), .Y(n3391) );
 NAND2X1TS U2610 ( .A(n3394), .A(n3394_n), .B(n3395), .B(n3395_n), .Y(n3393_n), .Y(n3393) );
 NAND2X1TS U2611 ( .A(n2714), .A(n2714_n), .B(n3396), .B(n3396_n), .Y(n3395_n), .Y(n3395) );
 NAND2X1TS U2612 ( .A(n2837), .A(n2837_n), .B(n2715), .B(n2715_n), .Y(n3396_n), .Y(n3396) );
 NAND2X1TS U2613 ( .A(n3560), .A(n3560_n), .B(n3561), .B(n3561_n), .Y(n2954_n), .Y(n2954) );
 NAND2X1TS U2614 ( .A(n2698), .A(n2698_n), .B(n3397), .B(n3397_n), .Y(n3394_n), .Y(n3394) );
 NAND2X1TS U2615 ( .A(n3398), .A(n3398_n), .B(n2772), .B(n2772_n), .Y(n3397_n), .Y(n3397) );
 NAND2X1TS U2616 ( .A(n3399), .A(n3399_n), .B(n3400), .B(n3400_n), .Y(n3392_n), .Y(n3392) );
 NAND2X1TS U2617 ( .A(n2725), .A(n2725_n), .B(n3401), .B(n3401_n), .Y(n3400_n), .Y(n3400) );
 NAND2X1TS U2618 ( .A(n2793), .A(n2793_n), .B(n2806), .B(n2806_n), .Y(n3401_n), .Y(n3401) );
 NAND2X1TS U2619 ( .A(n3408), .A(n3408_n), .B(n3409), .B(n3409_n), .Y(n3407_n), .Y(n3407) );
 NAND2X1TS U2620 ( .A(n2707), .A(n2707_n), .B(n3428), .B(n3428_n), .Y(n3096_n), .Y(n3096) );
 NAND2X1TS U2621 ( .A(n3414), .A(n3414_n), .B(n3415), .B(n3415_n), .Y(n3406_n), .Y(n3406) );
 NAND2X1TS U2622 ( .A(n2697), .A(n2697_n), .B(n2722), .B(n2722_n), .Y(n3288_n), .Y(n3288) );
 NAND2X1TS U2623 ( .A(n2899), .A(n2899_n), .B(n3586), .B(n3586_n), .Y(n3398_n), .Y(n3398) );
 NAND2X1TS U2624 ( .A(n2912), .A(n2912_n), .B(n2895), .B(n2895_n), .Y(n3527_n), .Y(n3527) );
 NAND2X1TS U2625 ( .A(n3422), .A(n3422_n), .B(n3423), .B(n3423_n), .Y(n3421_n), .Y(n3421) );
 NAND2X1TS U2626 ( .A(n2738), .A(n2738_n), .B(n3424), .B(n3424_n), .Y(n3423_n), .Y(n3423) );
 NAND2X1TS U2627 ( .A(n2801), .A(n2801_n), .B(n2719), .B(n2719_n), .Y(n3424_n), .Y(n3424) );
 NAND2X1TS U2628 ( .A(n2909), .A(n2909_n), .B(n2889), .B(n2889_n), .Y(n3524_n), .Y(n3524) );
 NAND2X1TS U2629 ( .A(n3555), .A(n3555_n), .B(n3459), .B(n3459_n), .Y(n3080_n), .Y(n3080) );
 NAND2X1TS U2630 ( .A(n2854), .A(n2854_n), .B(n3425), .B(n3425_n), .Y(n3422_n), .Y(n3422) );
 NAND2X1TS U2631 ( .A(n2801), .A(n2801_n), .B(n2780), .B(n2780_n), .Y(n3425_n), .Y(n3425) );
 NAND2X1TS U2632 ( .A(n2911), .A(n2911_n), .B(n3570), .B(n3570_n), .Y(n3569_n), .Y(n3569) );
 NAND2X1TS U2633 ( .A(n2893), .A(n2893_n), .B(n3428), .B(n3428_n), .Y(n3427_n), .Y(n3427) );
 MXI2X1TS U2634 ( .A(n3429), .A(n3429_n), .B(n2744), .B(n2744_n), .S0(n2905), .S0(n2905_n), .Y(n3426_n), .Y(n3426) );
 NAND2X1TS U2635 ( .A(n3560), .A(n3560_n), .B(n3587), .B(n3587_n), .Y(n2945_n), .Y(n2945) );
 NAND2X1TS U2636 ( .A(n2728), .A(n2728_n), .B(n2824), .B(n2824_n), .Y(n3429_n), .Y(n3429) );
 NAND2X1TS U2637 ( .A(n2895), .A(n2895_n), .B(n3562), .B(n3562_n), .Y(n3578_n), .Y(n3578) );
endmodule

